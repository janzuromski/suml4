�csklearn.ensemble._forest
RandomForestClassifier
q )�q}q(X   base_estimatorqcsklearn.tree._classes
DecisionTreeClassifier
q)�q}q(X	   criterionqX   giniqX   splitterq	X   bestq
X	   max_depthqNX   min_samples_splitqKX   min_samples_leafqKX   min_weight_fraction_leafqG        X   max_featuresqNX   max_leaf_nodesqNX   random_stateqNX   min_impurity_decreaseqG        X   class_weightqNX	   ccp_alphaqG        X   _sklearn_versionqX   1.0.2qubX   n_estimatorsqKX   estimator_paramsq(hhhhhhhhhhtqX	   bootstrapq�X	   oob_scoreq�X   n_jobsqNhNX   verboseqK X
   warm_startq�hNX   max_samplesqNhhhKhKhKhG        hX   autoq hNhG        hG        X   feature_names_in_q!cnumpy.core.multiarray
_reconstruct
q"cnumpy
ndarray
q#K �q$Cbq%�q&Rq'(KK�q(cnumpy
dtype
q)X   O8q*���q+Rq,(KX   |q-NNNJ����J����K?tq.b�]q/(X   Pclassq0X   Sexq1X   Ageq2X   SibSpq3X   Parchq4X   Fareq5X   Embarkedq6etq7bX   n_features_in_q8KX
   n_outputs_q9KX   classes_q:h"h#K �q;h%�q<Rq=(KK�q>h)X   i8q?���q@RqA(KX   <qBNNNJ����J����K tqCb�C               qDtqEbX
   n_classes_qFKX   base_estimator_qGhX   estimators_qH]qI(h)�qJ}qK(hhh	h
hKhKhKhG        hh hNhJ���*hG        hNhG        h8Kh9Kh:h"h#K �qLh%�qMRqN(KK�qOh)X   f8qP���qQRqR(KhBNNNJ����J����K tqSb�C              �?qTtqUbhFcnumpy.core.multiarray
scalar
qVhAC       qW�qXRqYX   max_features_qZKX   tree_q[csklearn.tree._tree
Tree
q\Kh"h#K �q]h%�q^Rq_(KK�q`hA�C       qatqbbK�qcRqd}qe(hKX
   node_countqfKcX   nodesqgh"h#K �qhh%�qiRqj(KKc�qkh)X   V56ql���qmRqn(Kh-N(X
   left_childqoX   right_childqpX   featureqqX	   thresholdqrX   impurityqsX   n_node_samplesqtX   weighted_n_node_samplesqutqv}qw(hoh)X   i8qx���qyRqz(KhBNNNJ����J����K tq{bK �q|hphzK�q}hqhzK�q~hrhRK�qhshRK �q�hthzK(�q�huhRK0�q�uK8KKtq�b�B�         *                 `f�$@���H.�?x           ��@       )                    @ҷ{�&�?�            �j@                           �?�@��u�?�            `j@                        �̌@���Q��?            �F@       
                    �?"pc�
�?            �@@                        �|�9@���}<S�?             7@������������������������       �                     @       	                    �?�t����?
             1@������������������������       �                      @������������������������       ��r����?	             .@                           �?���Q��?             $@                        ���@X�<ݚ�?             "@������������������������       �                      @������������������������       �և���X�?             @������������������������       �                     �?������������������������       �        	             (@                           �?���O1��?j            �d@                        P�J@     ��?             @@                           �? 	��p�?             =@                           �?�����H�?             2@������������������������       ��t����?             1@������������������������       �                     �?������������������������       �                     &@                        �|Y=@�q�q�?             @������������������������       �                     �?������������������������       �                      @       "                 �?�@�����?S            �`@                        ���@�8��8��?.             R@                            @�חF�P�?             ?@������������������������       �                     @������������������������       �z�G�z�?             9@        !                    �?��Y��]�?            �D@������������������������       �                     C@������������������������       ��q�q�?             @#       &                 0SE @j�g�y�?%             O@$       %                 ��) @�q�q�?             H@������������������������       ���Hg���?            �F@������������������������       �                     @'       (                   �;@@4և���?	             ,@������������������������       �                     (@������������������������       �      �?              @������������������������       �                     @+       J                    �?LGz���?�             x@,       7                    �?��&�?n            �f@-       2                   �H@HP�s��?              I@.       1                  S�-@���7�?             F@/       0                     @�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     C@3       6                    J@�q�q�?             @4       5                 ��Ca@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @8       C                    @d9q
$�?N            ``@9       @                 ���a@K�(i�?D            @]@:       =                    @��2(&�?A            �[@;       <                   `2@4��?�?>             Z@������������������������       ��GN�z�?             F@������������������������       �        %             N@>       ?                    @r�q��?             @������������������������       �                     @������������������������       �                     �?A       B                    <@և���X�?             @������������������������       �                     @������������������������       �                     @D       I                 ���d@����X�?
             ,@E       F                 ��T?@�C��2(�?	             &@������������������������       �                     @G       H                    %@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @K       X                    �?���?�            �i@L       U                    �?�X���?             F@M       R                     �?�4F����?            �D@N       O                   �8@d��0u��?             >@������������������������       �                     @P       Q                    �?r�q��?             8@������������������������       �                     *@������������������������       �                     &@S       T                   �;@"pc�
�?             &@������������������������       �                      @������������������������       �                     "@V       W                  "&d@�q�q�?             @������������������������       �                      @������������������������       �                     �?Y       b                    @��<b���?f             d@Z       _                 03�U@tk~X���?]             b@[       ^                    @\��I�h�?W             a@\       ]                     �?�F.< �?T            �`@������������������������       �p�v>��?            �G@������������������������       �z�G�z�?8            @U@������������������������       �                     @`       a                 03c@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �        	             1@q�tq�bX   valuesq�h"h#K �q�h%�q�Rq�(KKcKK�q�hR�B0       �u@     �o@      d@      K@      d@     �I@      2@      ;@      @      ;@       @      5@              @       @      .@               @       @      *@      @      @      @      @               @      @      @              �?      (@             �a@      8@      =@      @      ;@       @      0@       @      .@       @      �?              &@               @      �?              �?       @             @\@      5@     �P@      @      :@      @      @              4@      @      D@      �?      C@               @      �?     �G@      .@      A@      ,@      A@      &@              @      *@      �?      (@              �?      �?              @     �g@     �h@     �@@     �b@      @      G@       @      E@       @      @              @       @                      C@       @      @       @      �?       @                      �?              @      =@     �Y@      3@     �X@      .@     �W@      $@     �W@      $@      A@              N@      @      �?      @                      �?      @      @      @                      @      $@      @      $@      �?      @              @      �?              �?      @                      @     `c@      I@      =@      .@      <@      *@      3@      &@      @              *@      &@      *@                      &@      "@       @               @      "@              �?       @               @      �?             �_@     �A@     @[@     �A@     �Z@      ?@     @Y@      ?@     �@@      ,@      Q@      1@      @              @      @              @      @              1@        q�tq�bubhhubh)�q�}q�(hhh	h
hKhKhKhG        hh hNhJ��IShG        hNhG        h8Kh9Kh:h"h#K �q�h%�q�Rq�(KK�q�hR�C              �?q�tq�bhFhVhAC       q��q�Rq�hZKh[h\Kh"h#K �q�h%�q�Rq�(KK�q�hA�C       q�tq�bK�q�Rq�}q�(hKhfKShgh"h#K �q�h%�q�Rq�(KKS�q�hn�B(         L                    @>U���?�           ��@                          �0@�ˡ��A�?u           ؁@                          �A@nM`����?             G@                           @�'�=z��?            �@@       
                    #@��}*_��?             ;@       	                    �?؇���X�?
             ,@                            @�<ݚ�?             "@������������������������       �                      @������������������������       �����X�?             @������������������������       �                     @                           �?�n_Y�K�?	             *@                          �-@      �?             @������������������������       �                     �?������������������������       �                     @                           �?�<ݚ�?             "@������������������������       �      �?              @������������������������       �                     �?������������������������       �                     @                        ���`@$�q-�?             *@������������������������       �                     &@                        �(\�?      �?              @������������������������       �                     �?������������������������       �                     �?       5                    �?�������?W           h�@       &                    �?�p�*��?�            �w@                           �?8�A�0��?G            �[@                           �?$�q-�?            �C@                           2@�C��2(�?            �@@������������������������       �                     �?������������������������       �      �?             @@������������������������       �                     @        #                    �?��UV�?+            �Q@!       "                   �6@ДX��?)             Q@������������������������       �և���X�?             @������������������������       ���GEI_�?%            �N@$       %                    6@�q�q�?             @������������������������       �                      @������������������������       �                     �?'       .                    �?�r*��v�?�            �p@(       +                     @V�a�� �?)             M@)       *                     �?�FVQ&�?            �@@������������������������       �                     $@������������������������       ����}<S�?             7@,       -                    �?���Q��?             9@������������������������       �X�<ݚ�?             2@������������������������       �����X�?             @/       2                   �8@��ނ�b�?�            �j@0       1                 �1@lGts��?$            �K@������������������������       ��	j*D�?
             *@������������������������       ����N8�?             E@3       4                     �?�8",�?f            �c@������������������������       ��ʻ����?             A@������������������������       ����?N            �^@6       A                    �?��J~��?]             b@7       :                   �2@x!'ǯ�?/            �R@8       9                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @;       >                  S�-@0)RH'�?,            @Q@<       =                    �?      �?              @������������������������       ��q�q�?             @������������������������       �                      @?       @                    �?85�}C�?%            �N@������������������������       � ���J��?            �C@������������������������       �"pc�
�?             6@B       G                     �?�ˡ�5��?.            �Q@C       D                   �:@\X��t�?             7@������������������������       �                      @E       F                    �?�ՙ/�?             5@������������������������       �r�q��?             @������������������������       �z�G�z�?	             .@H       I                 �|�<@ �q�q�?              H@������������������������       �                     4@J       K                    @@@4և���?             <@������������������������       �8�Z$���?
             *@������������������������       �        	             .@M       R                    @ 	��p�?             =@N       O                 ��T?@����X�?             @������������������������       �                     @P       Q                 pf�C@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     6@q�tq�bh�h"h#K �q�h%�q�Rq�(KKSKK�q�hR�B0       @v@     �n@     �t@     @n@      1@      =@      0@      1@      $@      1@       @      (@       @      @               @       @      @              @       @      @      �?      @      �?                      @      @       @      @       @      �?              @              �?      (@              &@      �?      �?              �?      �?             �s@     �j@     �m@     �a@     @P@     �F@      @      B@      @      >@      �?               @      >@              @      O@      "@     �N@      @      @      @     �L@      @      �?       @               @      �?             �e@     @X@      (@      G@       @      ?@              $@       @      5@      $@      .@       @      $@       @      @      d@     �I@     �H@      @      "@      @      D@       @      \@     �F@      3@      .@     @W@      >@     �R@     �Q@      .@     �M@      @      �?              �?      @              &@      M@      @       @      @       @       @              @      L@      �?      C@      @      2@     �M@      (@      *@      $@               @      *@       @      �?      @      (@      @      G@       @      4@              :@       @      &@       @      .@              ;@       @      @       @      @              �?       @               @      �?              6@        q�tq�bubhhubh)�q�}q�(hhh	h
hKhKhKhG        hh hNhJu8�vhG        hNhG        h8Kh9Kh:h"h#K �q�h%�q�Rq�(KK�q�hR�C              �?q�tq�bhFhVhAC       q��q�Rq�hZKh[h\Kh"h#K �q�h%�q�Rq�(KK�q�hA�C       q�tq�bK�q�Rq�}q�(hKhfKwhgh"h#K �q�h%�q�Rq�(KKw�q�hn�B         2                    �?���ׁs�?n           ��@       #                    �?d�
��?K            �`@                           �?���@M^�?2            @W@                           �?\-��p�?             =@       
                     @HP�s��?             9@       	                     �?�nkK�?             7@                        �iE@�X�<ݺ?
             2@������������������������       �                     �?������������������������       �        	             1@������������������������       �                     @                        ��%@      �?              @������������������������       �                     �?������������������������       �                     �?                           �?      �?             @                          �>@      �?              @������������������������       �                     �?������������������������       �                     �?                        �|Y=@      �?              @������������������������       �                     �?������������������������       �                     �?                        ��UO@     8�?              P@                          @@      �?             L@������������������������       �                     ,@                            @r�q��?             E@                            �? ��WV�?             :@������������������������       ����N8�?	             5@������������������������       �                     @                        �|Y=@      �?             0@������������������������       �                     @������������������������       �                     $@                            �?      �?              @������������������������       �                     @!       "                 0wff@z�G�z�?             @������������������������       �                     @������������������������       �                     �?$       1                    �?�	j*D�?            �C@%       0                   �A@4�B��?            �B@&       +                    �?���Q��?             4@'       (                   �,@�q�q�?             .@������������������������       �                      @)       *                   �U@�θ�?	             *@������������������������       �ףp=
�?             $@������������������������       ��q�q�?             @,       /                 �|Y6@���Q��?             @-       .                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �        	             1@������������������������       �                      @3       d                     @����3��?#           @}@4       I                    �?�2�,��?~             i@5       B                   �;@�ݜ�?4            �S@6       ;                    �?��R[s�?            �A@7       :                    �?@4և���?	             ,@8       9                     �?؇���X�?             @������������������������       �                     @������������������������       ��q�q�?             @������������������������       �                     @<       ?                   �8@�ՙ/�?             5@=       >                 ���`@$�q-�?	             *@������������������������       �                     "@������������������������       �      �?             @@       A                    <@      �?              @������������������������       �                     @������������������������       ��q�q�?             @C       H                    �? qP��B�?            �E@D       E                    �?������?             B@������������������������       �                     @F       G                   �B@Pa�	�?            �@@������������������������       �                     7@������������������������       �ףp=
�?             $@������������������������       �                     @J       W                    �?03�Z*!�?J            �^@K       R                   �C@r�q��?:             X@L       O                   �?@؇>���?&            @P@M       N                   �;@��2(&�?             F@������������������������       ��X�<ݺ?             2@������������������������       ����B���?             :@P       Q                     �?�G��l��?
             5@������������������������       �����X�?             @������������������������       �X�Cc�?             ,@S       V                    �?�g�y��?             ?@T       U                   �=@���7�?             6@������������������������       �        
             0@������������������������       �r�q��?             @������������������������       �                     "@X       ]                    �?|��?���?             ;@Y       Z                    -@D�n�3�?             3@������������������������       �                     "@[       \                    �?z�G�z�?             $@������������������������       �                     @������������������������       ��q�q�?             @^       a                     �?      �?              @_       `                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?b       c                   `<@z�G�z�?             @������������������������       �                     @������������������������       �                     �?e       v                    @@�h�|5�?�            �p@f       m                  sW@
�cՔ��?�            @n@g       l                 ���@؇���X�?            �A@h       k                    ;@�d�����?
             3@i       j                   �5@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     (@������������������������       �                     0@n       u                    @��/�?            �i@o       r                    �?�q�q�?|             i@p       q                 X�lA@�P�*�?#             O@������������������������       ��F�j��?            �J@������������������������       �                     "@s       t                   �/@Ɔdq��?Y            `a@������������������������       ����"͏�?G            �[@������������������������       �      �?             <@������������������������       �                     @������������������������       �                     9@q�tq�bh�h"h#K �q�h%�q�Rq�(KKwKK�q�hR�Bp       �v@     @m@     @Q@     �O@     �L@      B@      @      9@       @      7@      �?      6@      �?      1@      �?                      1@              @      �?      �?              �?      �?               @       @      �?      �?              �?      �?              �?      �?              �?      �?             �J@      &@     �H@      @      ,@             �A@      @      9@      �?      4@      �?      @              $@      @              @      $@              @      @      @              �?      @              @      �?              (@      ;@      (@      9@      (@       @      $@      @               @      $@      @      "@      �?      �?       @       @      @       @      �?              �?       @                       @              1@               @     �r@     `e@     �Y@     �X@      $@      Q@      "@      :@      �?      *@      �?      @              @      �?       @              @       @      *@      �?      (@              "@      �?      @      @      �?      @               @      �?      �?      E@      �?     �A@              @      �?      @@              7@      �?      "@              @      W@      ?@     �S@      1@     �H@      0@      C@      @      1@      �?      5@      @      &@      $@       @      @      "@      @      >@      �?      5@      �?      0@              @      �?      "@              *@      ,@       @      &@              "@       @       @      @              @       @      @      @      �?       @               @      �?              @      �?      @                      �?     `h@      R@     @e@      R@      >@      @      ,@      @       @      @       @                      @      (@              0@             �a@     �P@     �`@     �P@      B@      :@      ;@      :@      "@             �X@     �D@      U@      ;@      ,@      ,@      @              9@        q�tq�bubhhubh)�q�}q�(hhh	h
hKhKhKhG        hh hNhJ�/GhG        hNhG        h8Kh9Kh:h"h#K �q�h%�q�Rq�(KK�q�hR�C              �?q�tq�bhFhVhAC       qՆq�Rq�hZKh[h\Kh"h#K �q�h%�q�Rq�(KK�q�hA�C       q�tq�bK�q�Rq�}q�(hKhfKUhgh"h#K �q�h%�q�Rq�(KKU�q�hn�B�                           `�X.@��gjN��?u           ��@                        ���+@�7���?�            �s@                        `f�$@v�u��?�            Pr@                           �?�%^�?�            �j@       
                 pF @>4և���?#             L@       	                    �?R���Q�?             D@                         s�@      �?             B@������������������������       �                     $@������������������������       �$��m��?             :@������������������������       �                     @                          #@      �?
             0@������������������������       �                      @                           �?      �?              @������������������������       �      �?             @������������������������       �                     @                           �?�S�%3��?j            �c@                            @$�Z����?c             c@������������������������       �                     @                         ��	@J�^y�?_             b@������������������������       �                     @������������������������       ���E�B��?^            �a@������������������������       �                     @                          �1@��Zy�?-            �S@������������������������       �                     &@                           �?�#}7��?'            �P@                        �J+@@i��M��?&            @P@                            @0�� ��?$            �O@������������������������       �¦	^_�?#             O@������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     3@!       :                     @�q���?�             r@"       -                    �?T+_Q���?z            �i@#       *                  "�b@ �#�Ѵ�?6            �U@$       )                    �?@	tbA@�?/            @Q@%       (                    �?`2U0*��?             9@&       '                    �?��S�ۿ?             .@������������������������       �؇���X�?             @������������������������       �                      @������������������������       �                     $@������������������������       �                     F@+       ,                    $@@�0�!��?             1@������������������������       �                     @������������������������       �                     ,@.       9                    @z�����?D            �]@/       4                     �?J�8���?C             ]@0       3                    �?t]����?2            �V@1       2                    �?      �?0             V@������������������������       �ҳ�wY;�?.            @U@������������������������       �                     @������������������������       �                     @5       6                    *@ �o_��?             9@������������������������       �                     @7       8                    �?ףp=
�?             4@������������������������       ��r����?
             .@������������������������       �                     @������������������������       �                     @;       F                 �̜3@j����?6            �T@<       =                    �?$��m��?             :@������������������������       �                     @>       A                    �?�\��N��?
             3@?       @                   @1@      �?              @������������������������       �                     @������������������������       �                     �?B       C                    �?���!pc�?             &@������������������������       �                     @D       E                    1@���Q��?             @������������������������       �                     @������������������������       �                      @G       N                    �?F�t�K��?'            �L@H       I                    ;@�eP*L��?             &@������������������������       �                     @J       K                    �?����X�?             @������������������������       �                     @L       M                    �?      �?             @������������������������       �                      @������������������������       �                      @O       P                    @�q��/��?             G@������������������������       �                      @Q       T                 ��p@@�?�'�@�?             C@R       S                    @��<b���?             7@������������������������       �                      @������������������������       �؇���X�?             5@������������������������       �        	             .@q�tq�bh�h"h#K �q�h%�q�Rq�(KKUKK�q�hR�BP       �v@     �m@     �k@     @V@     �i@     @V@      d@     �K@      7@     �@@      "@      ?@      "@      ;@              $@      "@      1@              @      ,@       @       @              @       @       @       @      @              a@      6@     @`@      6@      @             �^@      6@              @     �^@      2@      @              F@      A@              &@      F@      7@      F@      5@      F@      3@      F@      2@              �?               @               @      3@             @a@     �b@     �T@     �^@      @     �T@      �?      Q@      �?      8@      �?      ,@      �?      @               @              $@              F@      @      ,@      @                      ,@     �S@      D@      S@      D@      M@     �@@     �K@     �@@     �K@      >@              @      @              2@      @              @      2@       @      *@       @      @              @             �K@      <@      "@      1@              @      "@      $@      �?      @              @      �?               @      @      @               @      @              @       @              G@      &@      @      @              @      @       @      @               @       @               @       @             �D@      @       @             �@@      @      2@      @               @      2@      @      .@        q�tq�bubhhubh)�q�}q�(hhh	h
hKhKhKhG        hh hNhJ�vJhG        hNhG        h8Kh9Kh:h"h#K �q�h%�q�Rq�(KK�q�hR�C              �?q�tq�bhFhVhAC       q��q�Rq�hZKh[h\Kh"h#K �q�h%�q�Rq�(KK�q�hA�C       q�tq�bK�q�Rq�}r   (hKhfKWhgh"h#K �r  h%�r  Rr  (KKW�r  hn�B                              �?.�W����?s           ��@                           �?��}����?i            �c@                           �?�lO���?d             c@                        0Cd=@�?�P�a�?,             N@                            �?�'�`d�?            �@@                          �G@�q�q�?             @������������������������       �                     �?������������������������       �                      @	                           �?r�q��?             >@
                            @�θ�?	             *@������������������������       �                      @������������������������       ����!pc�?             &@                        �&�@�t����?             1@������������������������       �                     �?������������������������       �      �?             0@������������������������       �                     ;@                           @�㙢�c�?8             W@                           �?*c̕6�?5            �U@                        �|Y=@4�{Y���?2            �T@                           �?�X����?             6@������������������������       �      �?             4@������������������������       �                      @                        ���Q@Xny��?&            �N@������������������������       �l�b�G��?#            �L@������������������������       �      �?             @                           �?      �?             @������������������������       �                     �?                             @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @!       8                 `f�$@ز�h��?
           �{@"       7                    @xr����?i            @f@#       0                   @@@��/eA��?h             f@$       +                   �?@�-x�j�?R            `a@%       (                   �;@A5Xo�?N            ``@&       '                   �9@�Q��k�?0             T@������������������������       �pH����?)            �P@������������������������       ���
ц��?             *@)       *                 �|�=@���J��?            �I@������������������������       �                     G@������������������������       �z�G�z�?             @,       -                 P�@      �?              @������������������������       �                     �?.       /                 @3�@؇���X�?             @������������������������       �r�q��?             @������������������������       �                     �?1       2                      @P�Lt�<�?             C@������������������������       �                     @3       4                   @C@Pa�	�?            �@@������������������������       �        
             0@5       6                 �?�@�IєX�?             1@������������������������       �                     &@������������������������       �r�q��?             @������������������������       �                     �?9       V                  ޽j@�q�q�?�            �p@:       I                 `��R@^,IA4V�?�            p@;       B                    �?j���� �?�            �m@<       ?                    �?\������?@            @Z@=       >                   �<@"�W1��?.            �T@������������������������       �
j*D>�?             :@������������������������       � �Cc}�?              L@@       A                 03;@
;&����?             7@������������������������       �      �?             (@������������������������       �"pc�
�?             &@C       F                    �?���>���?Q            �`@D       E                     �?�㙢�c�?G            �\@������������������������       ��������?             A@������������������������       ��
��P�?1            @T@G       H                    @�����H�?
             2@������������������������       �                      @������������������������       �                     0@J       O                    �?p�ݯ��?             3@K       L                    �?؇���X�?             @������������������������       �                     @M       N                    5@      �?              @������������������������       �                     �?������������������������       �                     �?P       S                 03�a@      �?             (@Q       R                    �?����X�?             @������������������������       �                     @������������������������       �      �?             @T       U                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @r  tr  bh�h"h#K �r  h%�r  Rr	  (KKWKK�r
  hR�Bp       �x@      j@     �T@     �R@     �T@     @Q@      @     �J@      @      :@       @      �?              �?       @              @      9@      @      $@               @      @       @       @      .@      �?              �?      .@              ;@      S@      0@     �Q@      0@     @Q@      ,@      .@      @      .@      @               @      K@      @     �J@      @      �?      @       @       @      �?              �?       @      �?                       @      @                      @     Ps@     �`@     `c@      7@     `c@      6@     �]@      5@     @]@      ,@     �P@      *@      N@      @      @      @      I@      �?      G@              @      �?      �?      @              �?      �?      @      �?      @              �?     �B@      �?      @              @@      �?      0@              0@      �?      &@              @      �?              �?     @c@     �[@     `b@     �[@     �a@     �X@      =@      S@      1@     @P@      &@      .@      @      I@      (@      &@      @      "@      "@       @     �[@      6@     �W@      4@      9@      "@     �Q@      &@      0@       @               @      0@              @      (@      �?      @              @      �?      �?              �?      �?              @      @       @      @              @       @       @      @      �?      @                      �?      @        r  tr  bubhhubh)�r  }r  (hhh	h
hKhKhKhG        hh hNhJ�p�IhG        hNhG        h8Kh9Kh:h"h#K �r  h%�r  Rr  (KK�r  hR�C              �?r  tr  bhFhVhAC       r  �r  Rr  hZKh[h\Kh"h#K �r  h%�r  Rr  (KK�r  hA�C       r  tr  bK�r  Rr  }r   (hKhfK]hgh"h#K �r!  h%�r"  Rr#  (KK]�r$  hn�BX         N                    @      �?~           ��@       -                     @�ܞ6���?e           ��@                        �5L@�a�n��?�            �q@                            �?h0�����?{            @i@       
                   @B@T�iA�?(            �Q@                           �?���Q��?            �A@������������������������       �                      @       	                    �?|��?���?             ;@������������������������       �z�G�z�?             @������������������������       ��eP*L��?             6@                         �>@4�2%ޑ�?            �A@                           �?D�n�3�?             3@������������������������       ���.k���?             1@������������������������       �                      @������������������������       �                     0@                           2@d�
��?S            �`@������������������������       �        	             ,@                           �? ��X��?J            �]@                           �?r�q��?             (@������������������������       �      �?             @������������������������       �                      @                           �?      �?C            �Z@������������������������       �                     @������������������������       �D;����?A            �Y@                           �?l��
I��?4            @T@                        ���a@@9G��?            �H@������������������������       �                    �E@                           �?�q�q�?             @������������������������       �                     @������������������������       �                      @       &                    �?     ��?             @@        #                   �7@j���� �?             1@!       "                  D�U@�q�q�?             @������������������������       �                     @������������������������       ��q�q�?             @$       %                    �?���!pc�?             &@������������������������       �                     @������������������������       ����Q��?             @'       *                    �?z�G�z�?             .@(       )                 03�T@�8��8��?	             (@������������������������       �                      @������������������������       �      �?             @+       ,                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?.       A                    �?T�iA�?�            �q@/       <                   @B@&ջ�{��?4            @R@0       5                    @�ՙ/�?-            �O@1       4                    @؇���X�?             @2       3                    �?�q�q�?             @������������������������       �      �?              @������������������������       �                     �?������������������������       �                     @6       9                 �̌@>4և���?(             L@7       8                 ���@���B���?             :@������������������������       �                     @������������������������       ��GN�z�?             6@:       ;                    �?���Q��?             >@������������������������       ����Q��?             $@������������������������       ��z�G��?             4@=       @                    @z�G�z�?             $@>       ?                   �K@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     �?B       M                 �T�E@�_�/�?�            �i@C       H                    �?���x��?�            �i@D       G                    �?��s����?             5@E       F                    �?R���Q�?             4@������������������������       �@�0�!��?             1@������������������������       �                     @������������������������       �                     �?I       J                    )@�_�����?q             g@������������������������       �                      @K       L                    �?�h�ഭ�?p            �f@������������������������       �                     7@������������������������       �XT�z�q�?c            �c@������������������������       �                      @O       R                      @������?            �B@P       Q                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?S       \                 �|Y?@�IєX�?             A@T       U                    �?Pa�	�?            �@@������������������������       �        	             .@V       [                    @�X�<ݺ?             2@W       X                 ��T?@r�q��?             @������������������������       �                     @Y       Z                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     (@������������������������       �                     �?r%  tr&  bh�h"h#K �r'  h%�r(  Rr)  (KK]KK�r*  hR�B�       pw@      l@     `u@     �k@      `@     `c@      Z@     �X@     �D@      =@      ,@      5@               @      ,@      *@      @      �?      $@      (@      ;@       @      &@       @      "@       @       @              0@             �O@     @Q@              ,@     �O@     �K@      $@       @       @       @       @             �J@     �J@              @     �J@      I@      8@     �L@       @     �G@             �E@       @      @              @       @              6@      $@      $@      @       @      @              @       @      �?       @      @      @               @      @      (@      @      &@      �?       @              @      �?      �?       @               @      �?             �j@     �P@      @@     �D@      8@     �C@      �?      @      �?       @      �?      �?              �?              @      7@     �@@      @      5@              @      @      1@      2@      (@      @      @      ,@      @       @       @       @      �?       @                      �?              �?     �f@      9@     �f@      7@      1@      @      1@      @      ,@      @      @                      �?     �d@      3@               @     �d@      1@      7@             �a@      1@               @     �@@      @      �?       @               @      �?              @@       @      @@      �?      .@              1@      �?      @      �?      @               @      �?              �?       @              (@                      �?r+  tr,  bubhhubh)�r-  }r.  (hhh	h
hKhKhKhG        hh hNhJ�R�7hG        hNhG        h8Kh9Kh:h"h#K �r/  h%�r0  Rr1  (KK�r2  hR�C              �?r3  tr4  bhFhVhAC       r5  �r6  Rr7  hZKh[h\Kh"h#K �r8  h%�r9  Rr:  (KK�r;  hA�C       r<  tr=  bK�r>  Rr?  }r@  (hKhfKchgh"h#K �rA  h%�rB  RrC  (KKc�rD  hn�B�         4                    �?8C�N��?           ��@                        039@��Hg���?�             l@                           �?�T��5m�?T            �`@                        P�>,@z�G�z�?             �F@                            @�FVQ&�?            �@@������������������������       �                     @                        �|�9@ 	��p�?             =@������������������������       �                     $@	       
                 �&B@�KM�]�?             3@������������������������       �؇���X�?
             ,@������������������������       �                     @                           �?�q�q�?	             (@                          �#@���|���?             &@������������������������       �                      @                         S�2@�<ݚ�?             "@������������������������       �      �?              @������������������������       �                     �?������������������������       �                     �?                           @��9܂�?4            @V@                           �?|jq��?1            �T@                           �?�S���,�?0            @T@                           @�ՙ/�?&            �O@������������������������       ��-ῃ�?%            �N@������������������������       �                      @                          �9@X�<ݚ�?
             2@������������������������       �؇���X�?             @������������������������       �"pc�
�?             &@������������������������       �                      @                           @r�q��?             @������������������������       �                     @������������������������       �                     �?        1                    @$�q-�?@            �V@!       *                 `f~B@`��F:u�?<            �U@"       '                     @     ��?             @@#       $                   �G@��S�ۿ?             >@������������������������       �                     9@%       &                 ���;@���Q��?             @������������������������       �                     @������������������������       �                      @(       )                 ��p@@      �?              @������������������������       �                     �?������������������������       �                     �?+       ,                  "�b@ �Jj�G�?&            �K@������������������������       �                    �G@-       .                    �?      �?              @������������������������       �                     @/       0                 03c@z�G�z�?             @������������������������       �                     �?������������������������       �                     @2       3                    @      �?             @������������������������       �                     �?������������������������       �                     @5       N                    �?Tb�u �?�            pw@6       7                    )@xR�L::�?�            �q@������������������������       �                     @8       A                    �?���˰�?�            �q@9       @                 `��,@�����?-            �P@:       =                     @�L���?            �B@;       <                 X�l@@      �?              @������������������������       �                     �?������������������������       �                     �?>       ?                    �? >�֕�?            �A@������������������������       ���S�ۿ?             .@������������������������       �P���Q�?             4@������������������������       �                     >@B       I                    ?@�ˡ�5��?�            �j@C       F                   �3@��F���?T            �`@D       E                    &@ �o_��?             9@������������������������       �j���� �?             1@������������������������       �                      @G       H                 `fF:@h�WH��?F             [@������������������������       ���s��??            �W@������������������������       ���
ц��?             *@J       M                    �?�G�z.�?5             T@K       L                 �Y5@:���u��?2            @S@������������������������       �                     &@������������������������       ��j�'�=�?*            �P@������������������������       �                     @O       V                    @      �?2             V@P       S                    �?և���X�?             ,@Q       R                     @      �?              @������������������������       �                     @������������������������       �                     @T       U                    @�q�q�?             @������������������������       �                     @������������������������       �                      @W       `                   �L@��G���?+            �R@X       _                    @�ˡ�5��?)            �Q@Y       \                    �?z�G�z�?"             N@Z       [                     @�2����?            �K@������������������������       �������?             A@������������������������       ����N8�?
             5@]       ^                 �|�6@���Q��?             @������������������������       �                     �?������������������������       �      �?             @������������������������       �                     &@a       b                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?rE  trF  bh�h"h#K �rG  h%�rH  RrI  (KKcKK�rJ  hR�B0       �v@     �m@     �K@     @e@      H@     �U@      "@      B@       @      ?@              @       @      ;@              $@       @      1@       @      (@              @      @      @      @      @               @      @       @      @      �?              �?              �?     �C@      I@      A@     �H@      A@     �G@      8@     �C@      6@     �C@       @              $@       @      �?      @      "@       @               @      @      �?      @                      �?      @      U@      @     �T@      @      =@       @      <@              9@       @      @              @       @              �?      �?              �?      �?              �?      K@             �G@      �?      @              @      �?      @      �?                      @      @      �?              �?      @             0s@      Q@      n@      G@              @      n@     �C@      P@      @      A@      @      �?      �?              �?      �?             �@@       @      ,@      �?      3@      �?      >@              f@      B@      ]@      1@      2@      @      $@      @       @             �X@      $@     �V@      @      @      @     �N@      3@      M@      3@      &@             �G@      3@      @             �P@      6@      @       @      @      @              @      @               @      @              @       @              N@      ,@     �M@      (@      H@      (@      G@      "@      :@       @      4@      �?       @      @      �?              �?      @      &@              �?       @               @      �?        rK  trL  bubhhubh)�rM  }rN  (hhh	h
hKhKhKhG        hh hNhJh��UhG        hNhG        h8Kh9Kh:h"h#K �rO  h%�rP  RrQ  (KK�rR  hR�C              �?rS  trT  bhFhVhAC       rU  �rV  RrW  hZKh[h\Kh"h#K �rX  h%�rY  RrZ  (KK�r[  hA�C       r\  tr]  bK�r^  Rr_  }r`  (hKhfKohgh"h#K �ra  h%�rb  Rrc  (KKo�rd  hn�BH         "                   �1@���ׁs�?t           ��@       	                    �?���L��?6            �S@                           �?��s����?             5@                        ���0@������?	             1@                          �,@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     $@������������������������       �                     @
                           �?�\��N��?+            �L@                            @��
P��?            �A@������������������������       �                     @                           �?����"�?             =@                           '@�eP*L��?             &@������������������������       �                     @������������������������       �                     @                           @�E��ӭ�?             2@                            @      �?              @������������������������       ��q�q�?             @������������������������       �                      @                           �?ףp=
�?	             $@������������������������       �      �?              @������������������������       �                      @                           !@8�A�0��?             6@                        pf�C@ףp=
�?             $@������������������������       �                      @                           @      �?              @������������������������       �                     �?������������������������       �                     �?                           @�q�q�?	             (@������������������������       �                     @        !                 ���3@�����H�?             "@������������������������       �                     �?������������������������       �                      @#       F                    �?X�ym�?>           P�@$       3                     @��q���?t            `f@%       ,                   �H@X�?٥�?B            �Y@&       '                    �?F|/ߨ�?7            @T@������������������������       �                     F@(       +                    �?@-�_ .�?            �B@)       *                   �7@�FVQ&�?            �@@������������������������       �                     �?������������������������       �      �?             @@������������������������       �                     @-       2                   �I@��2(&�?             6@.       /                 03[;@�q�q�?             "@������������������������       �                     @0       1                 ��Ca@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     *@4       A                 м[8@:W��S��?2             S@5       <                 ��.@�ʻ����?.             Q@6       9                    �?(옄��?              G@7       8                 @3�@�\��N��?             C@������������������������       ���<b���?             7@������������������������       ��r����?
             .@:       ;                    �?      �?              @������������������������       �z�G�z�?             @������������������������       �                     @=       >                    5@�GN�z�?             6@������������������������       �                     @?       @                    C@�X�<ݺ?             2@������������������������       �                     1@������������������������       �                     �?B       C                 X��@@      �?              @������������������������       �                     @D       E                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?G       X                     �?|��Y���?�            pu@H       O                    �?�������?0            �V@I       J                   �8@4?,R��?             B@������������������������       �                      @K       L                    :@�>4և��?             <@������������������������       �                      @M       N                  �>@ȵHPS!�?             :@������������������������       �                     $@������������������������       �     ��?             0@P       W                    �?l��
I��?             K@Q       T                   @B@�#ʆA��?            �J@R       S                 �|�<@      �?             0@������������������������       �                      @������������������������       �և���X�?
             ,@U       V                    �?$G$n��?            �B@������������������������       �؇���X�?            �A@������������������������       �                      @������������������������       �                     �?Y       b                    �?pe7����?�            �o@Z       [                   @9@�θ�?             :@������������������������       �                     @\       _                 �̼*@�LQ�1	�?             7@]       ^                   @@�IєX�?             1@������������������������       ������H�?             "@������������������������       �                      @`       a                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @c       h                 �|�=@��)jO�?�            `l@d       g                    �?`�q�0ܴ?X            �a@e       f                    $@P#aE�?R            �`@������������������������       �t��ճC�?:             V@������������������������       �                    �F@������������������������       �                      @i       l                   @A@�4���L�?2            �U@j       k                    �?�ՙ/�?             5@������������������������       �      �?	             ,@������������������������       �؇���X�?             @m       n                    �?��ɉ�?&            @P@������������������������       �D>�Q�?             J@������������������������       �                     *@re  trf  bh�h"h#K �rg  h%�rh  Rri  (KKoKK�rj  hR�B�       �v@     @m@      ?@     �G@      @      1@      @      *@      @      @              @      @                      $@              @      ;@      >@      2@      1@              @      2@      &@      @      @      @                      @      *@      @      @      @       @      @       @              "@      �?      @      �?       @              "@      *@      �?      "@               @      �?      �?              �?      �?               @      @              @       @      �?              �?       @             �t@     `g@      E@      a@      @     �X@       @     �S@              F@       @     �A@       @      ?@      �?              �?      ?@              @      @      3@      @      @              @      @       @      @                       @              *@     �B@     �C@      >@      C@      9@      5@      2@      4@      @      2@      *@       @      @      �?      @      �?      @              @      1@      @              �?      1@              1@      �?              @      �?      @               @      �?       @                      �?     Pr@      I@     @Q@      5@      ?@      @       @              7@      @               @      7@      @      $@              *@      @      C@      0@      C@      .@      @      $@               @      @       @      @@      @      >@      @       @                      �?      l@      =@      4@      @              @      4@      @      0@      �?       @      �?       @              @       @               @      @             �i@      7@     �`@      @     �_@      @     �T@      @     �F@               @             @Q@      1@      *@       @      @      @      @      �?      L@      "@     �E@      "@      *@        rk  trl  bubhhubh)�rm  }rn  (hhh	h
hKhKhKhG        hh hNhJ�{�[hG        hNhG        h8Kh9Kh:h"h#K �ro  h%�rp  Rrq  (KK�rr  hR�C              �?rs  trt  bhFhVhAC       ru  �rv  Rrw  hZKh[h\Kh"h#K �rx  h%�ry  Rrz  (KK�r{  hA�C       r|  tr}  bK�r~  Rr  }r�  (hKhfKghgh"h#K �r�  h%�r�  Rr�  (KKg�r�  hn�B�         (                    �?X���[�?~           ��@       '                   @O@ �\��?o             d@                          �2@�J���?l            @c@                           �?������?             1@                        ج:#@8�Z$���?	             *@������������������������       �                     �?       
                    �?�8��8��?             (@       	                     @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @                          p2@      �?             @������������������������       �                      @������������������������       �                      @                           �?������?_             a@                            @և���X�?D            �X@                           �?      �?             @@������������������������       �        	             .@                           �?�IєX�?             1@������������������������       �                     &@������������������������       �r�q��?             @                           �?����e��?.            �P@                           �?���B���?             :@������������������������       ��q�q�?             8@������������������������       �                      @                          �+@      �?             D@������������������������       ���-�=��?            �C@������������������������       �                     �?       "                   @G@�e����?            �C@       !                   �C@      �?             >@                            �?���Q��?             9@������������������������       ��r����?
             .@������������������������       �z�G�z�?	             $@������������������������       �                     @#       $                    �?�����H�?             "@������������������������       �                     @%       &                   �H@r�q��?             @������������������������       �                     @������������������������       ��q�q�?             @������������������������       �                     @)       6                    @<��_�&�?           p{@*       1                    @z�G�z�?             4@+       0                    �?@4և���?	             ,@,       -                    �?r�q��?             @������������������������       �                     @.       /                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @2       3                    �?      �?             @������������������������       �                     �?4       5                 �̤=@���Q��?             @������������������������       �                      @������������������������       �                     @7       P                     @j��E�?           0z@8       G                   @E@�m����?m             f@9       @                    �?��R�?k�?S            �a@:       =                 03�a@�IєX�?%             Q@;       <                   �;@      �?"             P@������������������������       ����}<S�?             7@������������������������       �                    �D@>       ?                    �?      �?             @������������������������       �                     �?������������������������       ��q�q�?             @A       D                   pT@��oh���?.            @R@B       C                 `fF)@��X���?+            @Q@������������������������       �                     0@������������������������       ��c�����?            �J@E       F                    �?      �?             @������������������������       �                     �?������������������������       �                     @H       K                   �'@tk~X��?             B@I       J                    �?      �?             @������������������������       �                     @������������������������       �                     �?L       M                    �?      �?             @@������������������������       �                      @N       O                 `ff:@��S�ۿ?             >@������������������������       �                     &@������������������������       ��KM�]�?             3@Q       ^                    �?��8PTJ�?�            @n@R       Y                    �?�^���U�?#            �L@S       V                   �;@d�
��?             F@T       U                    �?�E��ӭ�?             2@������������������������       ��z�G��?             $@������������������������       �      �?              @W       X                   #@�	j*D�?             :@������������������������       �                     &@������������������������       ���S���?	             .@Z       [                    @$�q-�?	             *@������������������������       �                      @\       ]                 ���3@z�G�z�?             @������������������������       �                     �?������������������������       �                     @_       f                    �?t��eh��?r             g@`       c                    �?� U ��?i            �e@a       b                    ?@�~g�>�?[            �b@������������������������       ��LQ�1	�?D            �\@������������������������       �<ݚ)�?             B@d       e                  �'@��2(&�?             6@������������������������       �      �?             @������������������������       �                     0@������������������������       �        	             (@r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKgKK�r�  hR�Bp        w@      m@     �T@     �S@      S@     �S@      @      *@       @      &@      �?              �?      &@      �?      @              @      �?                       @       @       @               @       @              R@     @P@      L@      E@      0@      0@              .@      0@      �?      &@              @      �?      D@      :@      @      5@      @      3@               @     �A@      @     �A@      @              �?      0@      7@      .@      .@      $@      .@       @      *@       @       @      @              �?       @              @      �?      @              @      �?       @      @             �q@     @c@      @      0@      �?      *@      �?      @              @      �?       @      �?                       @               @      @      @      �?               @      @       @                      @     �q@     @a@     �V@     �U@     �N@      T@      @      P@       @      O@       @      5@             �D@       @       @              �?       @      �?     �L@      0@      L@      *@      0@              D@      *@      �?      @      �?                      @      =@      @      �?      @              @      �?              <@      @               @      <@       @      &@              1@       @     �g@     �I@     �A@      6@      7@      5@      @      *@      @      @       @      @      2@       @      &@              @       @      (@      �?       @              @      �?              �?      @             �c@      =@      b@      =@     @_@      :@      Y@      .@      9@      &@      3@      @      @      @      0@              (@        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hKhKhKhG        hh hNhJ2�8 hG        hNhG        h8Kh9Kh:h"h#K �r�  h%�r�  Rr�  (KK�r�  hR�C              �?r�  tr�  bhFhVhAC       r�  �r�  Rr�  hZKh[h\Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hA�C       r�  tr�  bK�r�  Rr�  }r�  (hKhfKihgh"h#K �r�  h%�r�  Rr�  (KKi�r�  hn�B�         2                    �?      �?�           ��@                          �2@ގ�H��?�            �x@                           $@>���Rp�?             =@                          �1@�eP*L��?             &@                           �?X�<ݚ�?             "@������������������������       �                      @       
                   �0@����X�?             @       	                 �̌!@      �?             @������������������������       ��q�q�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @                            �?�����H�?
             2@������������������������       �                     @                           �?"pc�
�?             &@                         S�(@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @       #                    �?�]<wr��?�            �v@       "                 `v�5@n�C���?C            �V@                           �?���|���?/            �P@                        ��	-@�S����?             3@                           �?�����H�?             2@������������������������       �                      @������������������������       �      �?
             0@������������������������       �                     �?                            @��V�I��?"            �G@                          �+@�t����?             1@������������������������       �"pc�
�?
             &@������������������������       �                     @        !                 �&B@d��0u��?             >@������������������������       ��<ݚ�?             "@������������������������       ���s����?             5@������������������������       �                     9@$       1                    �?�@�' �?�            0q@%       *                   �8@��2(&�?�            �p@&       '                    �?�}�+r��?"            �L@������������������������       �                     $@(       )                   �3@=QcG��?            �G@������������������������       �r�q��?             @������������������������       �������?            �D@+       .                    �?0)RH'�?y            �i@,       -                 �|Y=@ ��WV�?             J@������������������������       �                      @������������������������       �                     I@/       0                     �?z�G�z�?\            `c@������������������������       �l��
I��?             ;@������������������������       �     ��?J             `@������������������������       �                     &@3       J                    �?�p ��?�            �i@4       A                    �?�������?H            �Y@5       8                    @z�G�z�?5             T@6       7                 ��1V@      �?             @������������������������       �                      @������������������������       �                      @9       <                    .@�S����?3             S@:       ;                 xFT!@"pc�
�?             &@������������������������       �                      @������������������������       �                     "@=       >                     �?P�2E��?,            @P@������������������������       �                     ;@?       @                    �?�˹�m��?             C@������������������������       �l��\��?             A@������������������������       �                     @B       C                     @8�A�0��?             6@������������������������       �                     @D       E                 ���0@�E��ӭ�?             2@������������������������       �                     @F       G                    �?�r����?             .@������������������������       �                     �?H       I                    @@4և���?             ,@������������������������       �z�G�z�?             @������������������������       �        	             "@K       X                    �?ڲ�-���?B            �Y@L       S                 �TQK@X�<ݚ�?             2@M       N                    +@z�G�z�?             $@������������������������       �                     �?O       P                     @�����H�?             "@������������������������       �                      @Q       R                    �?؇���X�?             @������������������������       �                      @������������������������       �z�G�z�?             @T       W                    �?      �?              @U       V                 �U�X@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @Y       f                 03�U@z�G�z�?7            @U@Z       _                    �?r�q��?4            �S@[       \                     �?��(\���?             D@������������������������       �                     @]       ^                   �9@l��\��?             A@������������������������       �r�q��?             (@������������������������       ����7�?             6@`       c                     @�d�����?             C@a       b                    �?��
ц��?	             *@������������������������       ��eP*L��?             &@������������������������       �                      @d       e                    @H%u��?             9@������������������������       ����Q��?             @������������������������       �                     4@g       h                   �g@և���X�?             @������������������������       �                     @������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKiKK�r�  hR�B�       pw@      l@     �p@     @_@      @      6@      @      @      @      @               @      @       @       @       @      �?       @      �?              @                       @       @      0@              @       @      "@       @       @               @       @                      @     pp@     �Y@      8@     �P@      8@      E@      @      0@       @      0@               @       @      ,@      �?              5@      :@       @      .@       @      "@              @      3@      &@       @      @      1@      @              9@     �m@      B@     �l@      B@      K@      @      $@              F@      @      @      �?     �C@       @     �e@     �@@      I@       @               @      I@              _@      ?@      3@       @     @Z@      7@      &@             @Z@      Y@      ;@     �R@      ,@     �P@       @       @               @       @              (@      P@      "@       @               @      "@              @      O@              ;@      @     �A@      @      ?@              @      *@      "@              @      *@      @              @      *@       @              �?      *@      �?      @      �?      "@             �S@      9@      $@       @       @       @              �?       @      �?       @              @      �?       @              @      �?       @      @       @       @               @       @                      @      Q@      1@     @P@      *@     �B@      @      @              ?@      @      $@       @      5@      �?      <@      $@      @      @      @      @               @      6@      @       @      @      4@              @      @              @      @        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hKhKhKhG        hh hNhJ���'hG        hNhG        h8Kh9Kh:h"h#K �r�  h%�r�  Rr�  (KK�r�  hR�C              �?r�  tr�  bhFhVhAC       r�  �r�  Rr�  hZKh[h\Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hA�C       r�  tr�  bK�r�  Rr�  }r�  (hKhfKmhgh"h#K �r�  h%�r�  Rr�  (KKm�r�  hn�B�         F                  x#J@���H.�?�           ��@       #                    �?��)�7�?E           `@                          @B@.��|\�?l            �e@                        `f�$@�(�.Y��?_            `b@       
                   �3@�eP*L��?             F@       	                    �?؇���X�?             @                        �Y5@�q�q�?             @������������������������       �                     �?������������������������       �      �?              @������������������������       �                     @                        �̌@��+��?            �B@                           �?��}*_��?             ;@������������������������       �                     @������������������������       ��G��l��?             5@                        @3�@ףp=
�?             $@������������������������       ��q�q�?             @������������������������       �                     @                        `f�)@4A�,��?@            �Y@������������������������       �                     ,@                            @@�h�|5�?8            @V@                          �+@ףp=
�?             I@������������������������       �������?             .@������������������������       ���?^�k�?            �A@                        �|Y=@Hث3���?            �C@������������������������       ��d�����?             3@������������������������       �      �?             4@       "                    �?�q�����?             9@       !                 `v7<@և���X�?             5@                           �?p�ݯ��?
             3@������������������������       �                     @                            �?��S���?	             .@������������������������       �և���X�?             ,@������������������������       �                     �?������������������������       �                      @������������������������       �                     @$       9                    �?]����?�            �t@%       ,                  s�@֢�<���?�            �q@&       +                    �?�FVQ&�?+            �P@'       (                     @��S�ۿ?)             N@������������������������       �                     @)       *                   �8@,�+�C�?%            �K@������������������������       �                     4@������������������������       �(N:!���?            �A@������������������������       �                     @-       2                     @�t�i�?�            �k@.       1                   �B@:	��ʵ�?@            �V@/       0                 ��$:@|��"J�?9            @T@������������������������       ����c���?#             J@������������������������       �8^s]e�?             =@������������������������       �                     "@3       6                    �?��ׂ�?P            ``@4       5                 �|�=@��p��?K            @^@������������������������       ��㙢�c�?7             W@������������������������       �J�8���?             =@7       8                   �4@z�G�z�?             $@������������������������       �                     @������������������������       ��q�q�?             @:       ?                    @��V#�?            �E@;       <                     @����X�?
             ,@������������������������       �                      @=       >                     @�q�q�?             @������������������������       �                      @������������������������       �                     @@       E                     @\-��p�?             =@A       D                    �?"pc�
�?             6@B       C                     @�	j*D�?	             *@������������������������       �                     �?������������������������       �      �?             (@������������������������       �                     "@������������������������       �                     @G       d                 ���g@��O5���??            �X@H       Y                    E@b:�&���?6            �T@I       R                      @�^����?'            �M@J       Q                  ��T@�>����?"             K@K       N                  D:T@PN��T'�?             ;@L       M                    �?�8��8��?             8@������������������������       ��IєX�?             1@������������������������       �؇���X�?             @O       P                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     ;@S       X                    �?���Q��?             @T       U                    ;@�q�q�?             @������������������������       �                     �?V       W                    >@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @Z       ]                   �G@�q�q�?             8@[       \                    �?      �?             @������������������������       �                     @������������������������       �                     �?^       _                    �?      �?             4@������������������������       �                     &@`       c                    �?X�<ݚ�?             "@a       b                 @�pX@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @e       f                    5@��S���?	             .@������������������������       �                     @g       l                     @�q�q�?             (@h       k                    @X�<ݚ�?             "@i       j                 X�,@@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKmKK�r�  hR�B�       �u@     �o@     Pt@      f@     �L@     �\@      F@     �Y@      4@      8@      �?      @      �?       @              �?      �?      �?              @      3@      2@      $@      1@              @      $@      &@      "@      �?       @      �?      @              8@     �S@              ,@      8@     @P@      @     �F@      @      &@      �?      A@      3@      4@      ,@      @      @      .@      *@      (@      "@      (@      @      (@              @      @       @      @       @      �?               @              @             �p@      O@     �m@      H@      O@      @      L@      @      @             �I@      @      4@              ?@      @      @              f@      F@     �R@      0@     @P@      0@     �F@      @      4@      "@      "@             �Y@      <@     �W@      :@      S@      0@      3@      $@       @       @      @              �?       @      =@      ,@      @      $@               @      @       @               @      @              9@      @      2@      @      "@      @              �?      "@      @      "@              @              7@     �R@      .@      Q@      @      J@      @      I@      @      7@       @      6@      �?      0@      �?      @       @      �?              �?       @                      ;@      @       @      �?       @              �?      �?      �?      �?                      �?       @               @      0@      @      �?      @                      �?      @      .@              &@      @      @       @      @              @       @              @               @      @      @              @      @      @      @      @      @      @                      @       @                      @r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hKhKhKhG        hh hNhJ�%mthG        hNhG        h8Kh9Kh:h"h#K �r�  h%�r�  Rr�  (KK�r�  hR�C              �?r�  tr�  bhFhVhAC       r�  �r�  Rr�  hZKh[h\Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hA�C       r�  tr�  bK�r�  Rr�  }r�  (hKhfKchgh"h#K �r�  h%�r�  Rr�  (KKc�r�  hn�B�         .                     @f����?z           ��@                           �?.�����?�            �p@                           @�IєX�?N            �]@                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @                           6@���"�?L             ]@       	                    �?ףp=
�?             >@������������������������       �                     @
                           �?      �?             8@                          �2@R���Q�?             4@������������������������       ������H�?
             2@������������������������       �      �?              @������������������������       �                     @                           �? qP��B�?8            �U@                        03�<@ ��ʻ��?,             Q@                            �?      �?
             0@������������������������       ��q�q�?             @������������������������       �                     *@������������������������       �        "             J@                          �8@�X�<ݺ?             2@������������������������       �                     &@                           �?؇���X�?             @������������������������       �                     @������������������������       �      �?              @                          �1@BA�V�?[            �b@������������������������       �                     @       #                 ��D:@�q�q�?W             b@                            �?d1<+�C�?)            @R@������������������������       �                     @       "                    �?��hJ,�?&             Q@        !                    �?D|U��@�?%            �P@������������������������       �     ��?$             P@������������������������       �                     @������������������������       �                     �?$       )                    �?��M��?.            �Q@%       (                     �?H.�!���?              I@&       '                    �?�q�q��?             H@������������������������       �        	             0@������������������������       �     ��?             @@������������������������       �                      @*       -                   @I@և���X�?             5@+       ,                     @��.k���?             1@������������������������       �     ��?             0@������������������������       �                     �?������������������������       �                     @/       D                    �?�r��5�?�            �t@0       ;                  ��8@h0�����?D            @Y@1       8                    C@�,�٧��?:            �S@2       7                    @z�7�Z�?7            @R@3       4                    @ޚ)�?6             R@������������������������       �                     "@5       6                    �?p�EG/��?0            �O@������������������������       ��������?             A@������������������������       �П[;U��?             =@������������������������       �                     �?9       :                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @<       =                    �?���7�?
             6@������������������������       �                     @>       ?                    @��S�ۿ?             .@������������������������       �                     @@       C                     @ףp=
�?             $@A       B                 ��T?@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @E       J                 �� @��}���?�            �l@F       G                    6@���Q��?             $@������������������������       �                     @H       I                   �B@�q�q�?             @������������������������       �                     @������������������������       �                      @K       Z                    �?�t����?�            �k@L       S                    �?\-��p�?j            �e@M       P                   �6@HP�s��?             9@N       O                    5@      �?             @������������������������       �                     �?������������������������       ��q�q�?             @Q       R                 ���@���N8�?             5@������������������������       �                     @������������������������       �@4և���?
             ,@T       W                 �?�@�׆���?W            �b@U       V                    �?���;QU�?)            @R@������������������������       ��z�G��?             $@������������������������       ��i�y�?#            �O@X       Y                 �T)D@�A+K&:�?.             S@������������������������       �DE��2{�?-            �R@������������������������       �                     �?[       b                    @`�q�0ܴ?             �G@\       _                    �? �#�Ѵ�?            �E@]       ^                    �?�C��2(�?             &@������������������������       �                     @������������������������       �z�G�z�?             @`       a                    �?      �?             @@������������������������       �                     3@������������������������       �$�q-�?             *@������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKcKK�r�  hR�B0       `w@     @l@     @^@     `b@      @      \@       @      �?              �?       @              @     �[@      @      ;@              @      @      5@      @      1@       @      0@      �?      �?              @       @      U@      �?     �P@      �?      .@      �?       @              *@              J@      �?      1@              &@      �?      @              @      �?      �?     �\@     �A@              @     �\@      >@     �O@      $@      @              M@      $@     �L@      $@      K@      $@      @              �?             �I@      4@     �C@      &@     �B@      &@      0@              5@      &@       @              (@      "@       @      "@      @      "@      �?              @             �o@     �S@      J@     �H@      ?@      H@      :@     �G@      9@     �G@              "@      9@      C@      "@      9@      0@      *@      �?              @      �?              �?      @              5@      �?      @              ,@      �?      @              "@      �?       @      �?       @                      �?      @              i@      >@      @      @      @               @      @              @       @             `h@      :@     �b@      8@      7@       @      @      �?      �?               @      �?      4@      �?      @              *@      �?     �_@      6@      Q@      @      @      @     �N@       @     �M@      1@     �M@      0@              �?     �F@       @     �D@       @      $@      �?      @              @      �?      ?@      �?      3@              (@      �?      @        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hKhKhKhG        hh hNhJ�@�hG        hNhG        h8Kh9Kh:h"h#K �r�  h%�r�  Rr�  (KK�r�  hR�C              �?r�  tr�  bhFhVhAC       r�  �r�  Rr�  hZKh[h\Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hA�C       r�  tr�  bK�r�  Rr�  }r   (hKhfKahgh"h#K �r  h%�r  Rr  (KKa�r  hn�B8         ,                    �?f����?�           ��@                            @��ނ�b�?�            �j@                           �?H*C�|F�?R             `@                        03�<@��sK�z�?N            �^@       
                     �?ףp=
�?#             N@                          �G@      �?              @������������������������       �                     @       	                    �?      �?             @������������������������       �                      @������������������������       �                      @                           �?$�q-�?             J@������������������������       �                     @                          �B@Hm_!'1�?            �H@������������������������       �@-�_ .�?            �B@������������������������       �r�q��?             (@                         "�b@ ������?+            �O@������������������������       �        &            �L@                        03c@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @       '                    @��}E��?<            �T@                         ��.@�;�vv��?5            @R@                          �>@l`N���?'            �J@                           �?
;&����?#             G@                        �&�)@D�n�3�?             3@������������������������       �������?             .@������������������������       �                     @                           �?�5��?             ;@������������������������       �\X��t�?             7@������������������������       �      �?             @������������������������       �                     @!       &                    @�z�G��?             4@"       #                 03�1@�<ݚ�?             2@������������������������       �                     @$       %                 �I5@���|���?             &@������������������������       �z�G�z�?             @������������������������       �                     @������������������������       �                      @(       +                 ��T?@�z�G��?             $@)       *                 pfv2@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                      @-       D                    �?�蜹���?�            @x@.       9                    �?4և����?!             L@/       6                    �?؇���X�?             E@0       1                 ���@      �?             D@������������������������       �                     (@2       5                 p�i@@�>4և��?             <@3       4                   `=@�GN�z�?             6@������������������������       �R���Q�?             4@������������������������       �                      @������������������������       �                     @7       8                 03/O@      �?              @������������������������       �                     �?������������������������       �                     �?:       =                   �9@      �?	             ,@;       <                   �5@r�q��?             @������������������������       �                     �?������������������������       �                     @>       C                    �?      �?              @?       @                   �E@؇���X�?             @������������������������       �                     @A       B                   �H@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?E       P                    $@�1/z��?�            �t@F       K                    @      �?             4@G       H                    @�n_Y�K�?             *@������������������������       �                     @I       J                    �?�����H�?             "@������������������������       �                      @������������������������       �                     �?L       M                    !@����X�?             @������������������������       �                     @N       O                 ���9@      �?             @������������������������       �                      @������������������������       �                      @Q       X                   �A@���c���?�            �s@R       W                   @@@T�Jy&�?�             m@S       V                    �?�c�ve��?�            �j@T       U                   �?@�:pΈ��?x             i@������������������������       �°	~��?t             h@������������������������       �և���X�?             @������������������������       �                     .@������������������������       �        
             2@Y       `                    �?��t���?7            �S@Z       ]                 ��Q:@:�&���?6            �S@[       \                    �?�C��2(�?              F@������������������������       �                     @������������������������       ���-�=��?            �C@^       _                     �?�t����?             A@������������������������       ��q�q�?             >@������������������������       �                     @������������������������       �                     �?r  tr  bh�h"h#K �r  h%�r  Rr	  (KKaKK�r
  hR�B       `w@     @l@     �I@      d@      @     �^@      @      ]@      @      K@       @      @              @       @       @       @                       @      @      H@              @      @     �F@       @     �A@       @      $@      �?      O@             �L@      �?      @      �?                      @              @      F@     �C@     �B@      B@      ?@      6@      8@      6@       @      &@      @      &@      @              0@      &@      *@      $@      @      �?      @              @      ,@      @      ,@              @      @      @      @      �?              @       @              @      @      @      �?              �?      @                       @     0t@     @P@     �E@      *@      B@      @     �A@      @      (@              7@      @      1@      @      1@      @               @      @              �?      �?      �?                      �?      @      @      �?      @      �?                      @      @       @      @      �?      @               @      �?              �?       @                      �?     �q@      J@      $@      $@       @      @              @       @      �?       @                      �?       @      @              @       @       @               @       @             �p@      E@     �i@      <@     `g@      <@     �e@      <@      e@      9@      @      @      .@              2@             @P@      ,@      P@      ,@      D@      @      @             �A@      @      8@      $@      4@      $@      @              �?        r  tr  bubhhubh)�r  }r  (hhh	h
hKhKhKhG        hh hNhJ�i[hG        hNhG        h8Kh9Kh:h"h#K �r  h%�r  Rr  (KK�r  hR�C              �?r  tr  bhFhVhAC       r  �r  Rr  hZKh[h\Kh"h#K �r  h%�r  Rr  (KK�r  hA�C       r  tr  bK�r  Rr  }r   (hKhfKYhgh"h#K �r!  h%�r"  Rr#  (KKY�r$  hn�Bx         ,                    �?*;L]n�?q           ��@       !                 ��H@,i��?�            �j@                        0C�>@     ��?g             d@                            @tk~X���?\             b@                           �?�X�<ݺ?              K@       	                   �B@��(\���?             D@                           �?XB���?             =@������������������������       �                     @������������������������       ����7�?             6@
                           �?"pc�
�?             &@������������������������       �      �?              @������������������������       ������H�?             "@������������������������       �                     ,@                           @�L�lRT�?<            �V@                           7@NP�<��?7            �T@                         �}"@�n`���?             ?@������������������������       �        	             1@������������������������       �և���X�?             ,@                        ��.@�n_Y�K�?#             J@������������������������       ��'�=z��?            �@@������������������������       ��S����?             3@                           �?؇���X�?             @������������������������       �                     �?������������������������       �                     @                           �?      �?             0@������������������������       �                     @                           �?r�q��?             (@������������������������       �                     �?                            @�C��2(�?             &@                           @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@"       +                      @ ��WV�?"             J@#       $                    �?���J��?!            �I@������������������������       �                     :@%       &                    �?`2U0*��?             9@������������������������       �                     ,@'       (                 pf�\@�C��2(�?             &@������������������������       �                     "@)       *                     @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?-       @                 �?�@��3��?�            @x@.       ?                    �?lZ�?��?E            @]@/       <                    �?���}<S�?D            �\@0       5                    �?��<nd�?@            @[@1       2                 �|�:@      �?
             0@������������������������       �                     @3       4                 �|�=@�8��8��?             (@������������������������       �      �?              @������������������������       �                     @6       9                    �?��y� �?6            @W@7       8                  s�@�8��8��?	             (@������������������������       �                     @������������������������       �؇���X�?             @:       ;                   �;@ wVX(6�?-            @T@������������������������       �؇���X�?            �A@������������������������       ��nkK�?             G@=       >                 ��@r�q��?             @������������������������       �                     @������������������������       ��q�q�?             @������������������������       �                      @A       P                    @�)Y���?�            �p@B       C                    ,@���t�E�?�            �n@������������������������       �                     @D       I                 @3�@d��0u��?�             n@E       F                   �:@�q�q�?             @������������������������       �                     �?G       H                   �A@z�G�z�?             @������������������������       �                     �?������������������������       �      �?             @J       M                   �8@x�����?�            @m@K       L                    �?HP�s��?             I@������������������������       ������?             E@������������������������       �                      @N       O                    �?�5��
J�?q             g@������������������������       �&^�)b�?            �E@������������������������       ��*/�8V�?Y            �a@Q       X                 ���A@ �q�q�?             8@R       S                    �?ףp=
�?             $@������������������������       �                      @T       U                 �̤=@      �?              @������������������������       �                     @V       W                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     ,@r%  tr&  bh�h"h#K �r'  h%�r(  Rr)  (KKYKK�r*  hR�B�       �v@     `m@     �G@     �d@     �F@     �\@     �A@     @[@      @     �I@      @     �B@      �?      <@              @      �?      5@       @      "@      �?      �?      �?       @              ,@      @@      M@      :@     �L@      @      9@              1@      @       @      4@      @@      1@      0@      @      0@      @      �?              �?      @              $@      @              @      $@       @              �?      $@      �?      �?      �?      �?                      �?      "@               @      I@      �?      I@              :@      �?      8@              ,@      �?      $@              "@      �?      �?      �?                      �?      �?             �s@     �Q@     �Z@      $@     @Z@      $@      Y@      "@      .@      �?      @              &@      �?      @      �?      @             @U@       @      &@      �?      @              @      �?     �R@      @      >@      @      F@       @      @      �?      @               @      �?       @             `j@      N@     �g@     �M@              @     �g@      J@       @      @      �?              �?      @              �?      �?      @     @g@      H@      G@      @      C@      @       @             �a@      F@     �A@       @     @Z@      B@      7@      �?      "@      �?       @              @      �?      @               @      �?              �?       @              ,@        r+  tr,  bubhhubh)�r-  }r.  (hhh	h
hKhKhKhG        hh hNhJ�ܱLhG        hNhG        h8Kh9Kh:h"h#K �r/  h%�r0  Rr1  (KK�r2  hR�C              �?r3  tr4  bhFhVhAC       r5  �r6  Rr7  hZKh[h\Kh"h#K �r8  h%�r9  Rr:  (KK�r;  hA�C       r<  tr=  bK�r>  Rr?  }r@  (hKhfKyhgh"h#K �rA  h%�rB  RrC  (KKy�rD  hn�Bx         2                    �?�T���N�?p           ��@       !                 03�S@�eT+��?�            0y@                           +@t��:���?�            �w@                        `f7@ףp=
�?             $@������������������������       �                     @                        0339@      �?             @������������������������       �                     �?������������������������       �                     @	                           �?���V��?�            �v@
                        pff@V8Ɓ���?�            0u@                        03�@�C��2(�?$            �K@������������������������       �                     4@                           �?؇���X�?            �A@������������������������       �������?             .@������������������������       �P���Q�?             4@                           �?�O����?�            �q@                          @,@؀�:M�?*            �R@������������������������       �      �?             E@������������������������       �     ��?             @@                           �?���L��?�            @j@������������������������       �      �?             B@������������������������       �&y�X���?n            �e@                        `v�5@և���X�?             <@                            @d}h���?	             ,@������������������������       �                      @                        �|Y=@�8��8��?             (@������������������������       ��q�q�?             @������������������������       �                     "@                            E@X�Cc�?             ,@                            �?ףp=
�?             $@������������������������       �      �?              @������������������������       �                      @������������������������       �                     @"       )                  ޅg@8�Z$���?             :@#       (                    �?�}�+r��?             3@$       '                 �|�9@$�q-�?             *@%       &                  D�[@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@������������������������       �                     @*       1                    �?և���X�?             @+       .                    �?�q�q�?             @,       -                    �?      �?             @������������������������       �                     @������������������������       �                     �?/       0                   �B@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?3       V                 м�9@P��mu��?u            �h@4       C                    �?H�U?B�?2            �T@5       :                    �?)O���?             B@6       9                  S�-@����X�?             @7       8                 �&�)@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @;       B                    @l��[B��?             =@<       ?                    �?
j*D>�?             :@=       >                    �?j���� �?
             1@������������������������       ����Q��?             .@������������������������       �      �?              @@       A                     @�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     @D       O                    �?��<b���?             G@E       J                    �?@�0�!��?             A@F       I                 �&�)@��s����?             5@G       H                 ��@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �        	             (@K       N                    �?8�Z$���?             *@L       M                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@P       Q                     @�q�q�?             (@������������������������       �                     �?R       S                 ��'@���|���?             &@������������������������       �                     @T       U                 �|Y?@և���X�?             @������������������������       �                     @������������������������       �                     @W       p                    @�LQ�1	�?C            �\@X       a                    �?J����?:            �X@Y       \                   �@@��a�n`�?             ?@Z       [                    �?"pc�
�?             &@������������������������       �                     "@������������������������       �                      @]       ^                 @�pX@P���Q�?             4@������������������������       �        
             0@_       `                    �?      �?             @������������������������       �                     @������������������������       �                     �?b       i                 03�;@.Lj���?'             Q@c       f                    �?8�Z$���?             :@d       e                    :@�X�<ݺ?	             2@������������������������       ��8��8��?             (@������������������������       �                     @g       h                    �?      �?              @������������������������       ����Q��?             @������������������������       �                     @j       m                    �?��6���?             E@k       l                     @�㙢�c�?             7@������������������������       �        
             3@������������������������       �                     @n       o                    @���y4F�?             3@������������������������       �                     @������������������������       �      �?             0@q       r                    �?      �?	             0@������������������������       �                     @s       t                 ��T?@z�G�z�?             $@������������������������       �                     @u       x                    @�q�q�?             @v       w                    @���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?rE  trF  bh�h"h#K �rG  h%�rH  RrI  (KKyKK�rJ  hR�B�       w@     �l@     @q@     �_@      q@     @Z@      �?      "@              @      �?      @      �?                      @     �p@      X@     �o@      U@      I@      @      4@              >@      @      &@      @      3@      �?     �i@     �S@      G@      <@      5@      5@      9@      @     �c@     �I@      2@      2@     �a@     �@@      0@      (@      &@      @               @      &@      �?       @      �?      "@              @      "@      �?      "@      �?      @               @      @              @      6@      �?      2@      �?      (@      �?      �?              �?      �?                      &@              @      @      @       @      @      �?      @              @      �?              �?      �?      �?                      �?      �?             @W@      Z@     �J@      =@      1@      3@       @      @       @       @               @       @                      @      .@      ,@      .@      &@      @      $@      @      "@      �?      �?       @      �?       @                      �?              @      B@      $@      <@      @      1@      @      @      @      @                      @      (@              &@       @      �?       @      �?                       @      $@               @      @      �?              @      @      @              @      @              @      @              D@     �R@      :@     @R@      @      <@       @      "@              "@       @              �?      3@              0@      �?      @              @      �?              7@     �F@      @      6@      �?      1@      �?      &@              @      @      @      @       @              @      3@      7@      @      3@              3@      @              .@      @              @      .@      �?      ,@       @      @               @       @      @              @       @      @       @               @      @              �?        rK  trL  bubhhubh)�rM  }rN  (hhh	h
hKhKhKhG        hh hNhJ��ThG        hNhG        h8Kh9Kh:h"h#K �rO  h%�rP  RrQ  (KK�rR  hR�C              �?rS  trT  bhFhVhAC       rU  �rV  RrW  hZKh[h\Kh"h#K �rX  h%�rY  RrZ  (KK�r[  hA�C       r\  tr]  bK�r^  Rr_  }r`  (hKhfKGhgh"h#K �ra  h%�rb  Rrc  (KKG�rd  hn�B�         (                   �'@���Q��?m           ��@                           �?�?a/��?�             o@                        `f�$@:2vz�M�?&            �N@                           �?\�����?!            �K@       
                 �|�=@��k��?            �J@       	                 @3�@�(�Tw��?            �C@                           .@@�0�!��?             A@������������������������       �                     �?������������������������       �6YE�t�?            �@@������������������������       �                     @                          #@@4և���?             ,@������������������������       �                     (@                           I@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @                           +@ .2��A�?q            �g@������������������������       �                     �?                        ��@x�kE�?p            `g@                            @�}��L�?)            �R@������������������������       �                     @                           �? ��ʻ��?&             Q@                        �|�9@P���Q�?
             4@������������������������       �                     @������������������������       �      �?             0@������������������������       �                     H@       !                 ��L@>4և�z�?G             \@                           4@�q�q�?             (@������������������������       �                      @                            �?�z�G��?             $@������������������������       �      �?             @������������������������       �                     @"       %                   �E@ףp=
�?@             Y@#       $                    �?DE�SA_�?=            @X@������������������������       ����}<S�?;             W@������������������������       �                     @&       '                 @3�@�q�q�?             @������������������������       �                     �?������������������������       �      �?              @)       F                    P@L�5���?�            �u@*       A                    @vZoz��?�            �u@+       :                     @0R>�x�?�            `t@,       3                    �?�R�G�?�            @o@-       0                   �J@2ox��?Z            �c@.       /                    �?�2��P��?B            �\@������������������������       �X&$�E�?7            �X@������������������������       �     ��?             0@1       2                   �6@���N8�?             E@������������������������       �      �?              @������������������������       �@�0�!��?             A@4       7                    �?~��|��?6            @W@5       6                    @�h����?              L@������������������������       �      �?              @������������������������       � 7���B�?             K@8       9                   �B@��+��?            �B@������������������������       ��q�q�?	             .@������������������������       �8�A�0��?             6@;       <                   �*@\�Uo��?4             S@������������������������       �                     @=       >                    #@*O���?2             R@������������������������       �                     &@?       @                   �6@�jTM��?+            �N@������������������������       �                     *@������������������������       �     ��?$             H@B       C                    �?�����?             5@������������������������       �                     �?D       E                 ���d@P���Q�?             4@������������������������       �                     3@������������������������       �                     �?������������������������       �                     @re  trf  bh�h"h#K �rg  h%�rh  Rri  (KKGKK�rj  hR�Bp       �v@      n@     `h@      K@      :@     �A@      :@      =@      8@      =@      &@      <@      @      <@      �?              @      <@      @              *@      �?      (@              �?      �?      �?                      �?       @                      @      e@      3@              �?      e@      2@     �R@      �?      @             �P@      �?      3@      �?      @              .@      �?      H@             �W@      1@      @      @       @              @      @      @      @              @     �V@      $@     @V@       @      U@       @      @              �?       @              �?      �?      �?     �d@     @g@      d@     @g@     �a@      g@      X@     @c@     �R@     �T@      P@     �I@     �N@      C@      @      *@      $@      @@      @      @      @      <@      6@     �Q@      @     �J@      �?      �?       @      J@      3@      2@      $@      @      "@      *@      G@      >@              @      G@      :@              &@      G@      .@      *@             �@@      .@      3@       @              �?      3@      �?      3@                      �?      @        rk  trl  bubhhubh)�rm  }rn  (hhh	h
hKhKhKhG        hh hNhJ�I�BhG        hNhG        h8Kh9Kh:h"h#K �ro  h%�rp  Rrq  (KK�rr  hR�C              �?rs  trt  bhFhVhAC       ru  �rv  Rrw  hZKh[h\Kh"h#K �rx  h%�ry  Rrz  (KK�r{  hA�C       r|  tr}  bK�r~  Rr  }r�  (hKhfKqhgh"h#K �r�  h%�r�  Rr�  (KKq�r�  hn�B�         6                 ��K.@�T���N�?�           ��@                           �?浛��t�?�            ps@                        @1,@^�JB=�?5            @T@                           �?�z�G��?-            �Q@       
                 `fV$@R=6�z�?+            @P@       	                 �|�=@��J�fj�?            �B@                           �?     ��?             @@������������������������       �R���Q�?             4@������������������������       ��q�q�?
             (@������������������������       �                     @                           �? �Cc}�?             <@                           �?H%u��?             9@������������������������       �                     @������������������������       �r�q��?             2@������������������������       �                     @                           1@���Q��?             @������������������������       �                     @������������������������       �                      @                            @�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@                        ��@�LQ�1	�?�            �l@                        �Y�@H�!b	�?2            @T@                            @�����?             E@������������������������       �                     "@                        �|�=@<���D�?            �@@                           �?�㙢�c�?             7@������������������������       �z�G�z�?
             .@������������������������       �      �?              @������������������������       �                     $@������������������������       �                    �C@        '                    �?��H�&p�?a            �b@!       &                 �R,@      �?
             4@"       #                 �|Y=@�t����?             1@������������������������       �                     @$       %                 �|Y?@؇���X�?             ,@������������������������       �z�G�z�?             $@������������������������       �                     @������������������������       �                     @(       /                 �Yu@�T|n�q�?W             `@)       ,                 �?$@��
ц��?	             *@*       +                 �|Y9@�q�q�?             @������������������������       �                     �?������������������������       �                      @-       .                 �|�>@���Q��?             $@������������������������       �      �?              @������������������������       �                      @0       3                   �D@X�
����?N             ]@1       2                    �? i���t�?B            �X@������������������������       ��KM�]�?@            �W@������������������������       �                     @4       5                   @G@�E��ӭ�?             2@������������������������       ��q�q�?             @������������������������       ��8��8��?             (@7       ^                     @�^3�l��?�            r@8       K                 ��gS@�d�K���?�             i@9       >                    �?vA����?[            ``@:       =                   �;@����?�?             �F@;       <                   �9@      �?             0@������������������������       �                     .@������������������������       �                     �?������������������������       �                     =@?       F                     �?^����?;            �U@@       C                    �?������?&            �I@A       B                    �?>��C��?             �E@������������������������       �"pc�
�?	             &@������������������������       �      �?             @@D       E                 `��Q@      �?              @������������������������       ����Q��?             @������������������������       �                     @G       H                    *@^������?            �A@������������������������       �                     &@I       J                    �? �q�q�?             8@������������������������       �                     "@������������������������       ���S�ۿ?             .@L       Y                    �?��R[s�?)            �Q@M       R                 �|�<@�'N��?#            �N@N       O                    �?      �?
             2@������������������������       �                     @P       Q                 �U�X@"pc�
�?             &@������������������������       ����Q��?             @������������������������       �                     @S       V                 ���b@&^�)b�?            �E@T       U                 ��)[@�?�'�@�?             C@������������������������       �z�G�z�?             9@������������������������       �        	             *@W       X                    �?���Q��?             @������������������������       �      �?             @������������������������       �                     �?Z       ]                    �?�����H�?             "@[       \                    6@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @_       j                    �?�0�~�4�?8             V@`       a                    9@X�Emq�?             �J@������������������������       �                     &@b       i                   @C@��6���?             E@c       f                 ���;@)O���?             B@d       e                    �?և���X�?             <@������������������������       �p�ݯ��?             3@������������������������       �X�<ݚ�?             "@g       h                    �?      �?              @������������������������       �r�q��?             @������������������������       �                      @������������������������       �                     @k       p                 03�7@��?^�k�?            �A@l       m                 �|�7@      �?              @������������������������       �                     @n       o                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     ;@r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKqKK�r�  hR�B       w@     �l@     �l@      T@      ?@      I@      5@     �H@      3@      G@      0@      5@      &@      5@      @      1@       @      @      @              @      9@      @      6@              @      @      .@              @       @      @              @       @              $@      �?              �?      $@              i@      >@     @S@      @      C@      @      "@              =@      @      3@      @      (@      @      @      �?      $@             �C@             �^@      :@      .@      @      (@      @              @      (@       @       @       @      @              @              [@      5@      @      @      �?       @      �?                       @      @      @      @       @               @     @Y@      .@      V@      $@     @U@      $@      @              *@      @       @      @      &@      �?     @a@     �b@     @T@      ^@     �O@      Q@      �?      F@      �?      .@              .@      �?                      =@      O@      8@     �C@      (@     �@@      $@      "@       @      8@       @      @       @      @       @      @              7@      (@              &@      7@      �?      "@              ,@      �?      2@      J@      1@      F@      "@      "@              @      "@       @      @       @      @               @     �A@      @     �@@      @      4@              *@      @       @       @       @      �?              �?       @      �?       @               @      �?                      @     �L@      ?@      7@      >@              &@      7@      3@      1@      3@      0@      (@      (@      @      @      @      �?      @      �?      @               @      @              A@      �?      @      �?      @               @      �?       @                      �?      ;@        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hKhKhKhG        hh hNhJ�5ShG        hNhG        h8Kh9Kh:h"h#K �r�  h%�r�  Rr�  (KK�r�  hR�C              �?r�  tr�  bhFhVhAC       r�  �r�  Rr�  hZKh[h\Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hA�C       r�  tr�  bK�r�  Rr�  }r�  (hKhfKYhgh"h#K �r�  h%�r�  Rr�  (KKY�r�  hn�Bx         6                     @����fg�?�           ��@                          �8@���6��?�            �p@                          �1@d��0u��?'             N@������������������������       �                     1@                           �?�^�����?            �E@                           �?� �	��?             9@       
                   �3@�8��8��?             (@       	                   �'@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@                            �?�θ�?	             *@������������������������       �                     @                           �?�z�G��?             $@������������������������       ��q�q�?             "@������������������������       �                     �?                           �?�����H�?             2@                            �?�<ݚ�?             "@                          �7@�q�q�?             @������������������������       �                      @������������������������       �                     �?                          p@@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@       +                  D<Q@r�h����?�            �i@       *                    �?�z�Ga�?`             d@       #                    �?��EidD�?_            �c@                            �?      �?             <@                          �G@"pc�
�?             &@������������������������       �                      @������������������������       ��q�q�?             @!       "                  �>@�t����?             1@������������������������       �ףp=
�?             $@������������������������       �և���X�?             @$       '                   �@@�[�}r�?L            ``@%       &                    :@�q�q�?>             [@������������������������       �$��m��?0            �S@������������������������       ����Q��?             >@(       )                    �?���}<S�?             7@������������������������       �                     ,@������������������������       ��<ݚ�?             "@������������������������       �                     �?,       5                   �O@��|�5��?#            �G@-       4                    �?"pc�
�?"             F@.       1                    �?�T|n�q�?!            �E@/       0                    �?4?,R��?             B@������������������������       �                     <@������������������������       �      �?              @2       3                    �?����X�?             @������������������������       �                     @������������������������       ��q�q�?             @������������������������       �                     �?������������������������       �                     @7       X                  ��8@+F�	��?�            �t@8       K                 P��%@�;ĝ6�?�            �q@9       B                 pF @�G�5��?�            �i@:       A                   @F@�>�p���?e             b@;       >                    �?���ʻ��?^             a@<       =                    �?���@��?            �B@������������������������       �4�2%ޑ�?            �A@������������������������       �                      @?       @                    �?����!�?D            �X@������������������������       �4\�����?=            @V@������������������������       �                     $@������������������������       �                     "@C       J                    �?��� ��?-             O@D       G                    �?\-��p�?*             M@E       F                   p"@ףp=
�?             $@������������������������       �                     @������������������������       ��q�q�?             @H       I                 ���"@8��8���?#             H@������������������������       �X�EQ]N�?             �E@������������������������       ����Q��?             @������������������������       �                     @L       Q                    �?R�����?.             T@M       P                 033.@�����?
             3@N       O                 �&�)@�q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     $@R       S                   �*@�u���?$            �N@������������������������       �                     @T       W                   �?@J��D��?!             K@U       V                    �?v�2t5�?            �D@������������������������       ��q�q�?             @������������������������       �\�Uo��?             C@������������������������       �                     *@������������������������       �                     G@r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKYKK�r�  hR�B�       �v@      m@     �^@      b@      *@     �G@              1@      *@      >@      &@      ,@      �?      &@      �?      �?              �?      �?                      $@      $@      @      @              @      @      @      @      �?               @      0@       @      @      �?       @               @      �?              �?      @              @      �?                      "@     @[@     �X@     �X@      O@     �X@     �N@      ,@      ,@       @      "@               @       @      �?      (@      @      "@      �?      @      @      U@     �G@     �O@     �F@     �I@      ;@      (@      2@      5@       @      ,@              @       @              �?      &@      B@       @      B@      @      B@      @      ?@              <@      @      @       @      @              @       @      �?      �?              @             �n@      V@     �h@      V@     �c@     �I@     �Y@     �E@     @W@     �E@       @      =@       @      ;@               @     @U@      ,@     �R@      ,@      $@              "@              K@       @      I@       @      "@      �?      @               @      �?     �D@      @      C@      @      @       @      @             �E@     �B@      @      *@      @      @              @      @                      $@     �B@      8@              @     �B@      1@      8@      1@      �?       @      7@      .@      *@              G@        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hKhKhKhG        hh hNhJ��HhG        hNhG        h8Kh9Kh:h"h#K �r�  h%�r�  Rr�  (KK�r�  hR�C              �?r�  tr�  bhFhVhAC       r�  �r�  Rr�  hZKh[h\Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hA�C       r�  tr�  bK�r�  Rr�  }r�  (hKhfKqhgh"h#K �r�  h%�r�  Rr�  (KKq�r�  hn�B�         6                    �?��H�}�?�           ��@                            @���BK�?�            �j@                           :@ (��?D            @\@                           �?(L���?            �E@                           �?�8��8��?             B@������������������������       �                     @       
                   �+@ףp=
�?             >@       	                    B@d}h���?             ,@������������������������       ��C��2(�?             &@������������������������       ��q�q�?             @������������������������       �        	             0@                           �?և���X�?             @                          �7@���Q��?             @������������������������       �                      @������������������������       �                     @                           ,@      �?              @������������������������       �                     �?������������������������       �                     �?                           �?`����֜?*            �Q@������������������������       �                     <@                           �?�Ń��̧?             E@������������������������       �                     >@                          �8@�8��8��?             (@������������������������       �                     &@������������������������       �                     �?       3                    @      �?C             Y@       *                 �|�=@|jq��?9            �T@       #                 @3�@<=�,S��?/            �Q@                         �|Y<@�C��2(�?            �@@                        �Y5@���7�?
             6@������������������������       �ףp=
�?             $@������������������������       �                     (@!       "                 �&B@"pc�
�?
             &@������������������������       �      �?              @������������������������       �                     @$       '                 ���.@؀�:M�?            �B@%       &                 P��%@�KM�]�?             3@������������������������       �                     *@������������������������       ��q�q�?             @(       )                    �?�q�q�?             2@������������������������       �ףp=
�?             $@������������������������       �      �?              @+       0                    �?�n_Y�K�?
             *@,       -                   @"@և���X�?             @������������������������       �                      @.       /                    J@z�G�z�?             @������������������������       �      �?              @������������������������       �                     @1       2                 �̤=@r�q��?             @������������������������       �                     @������������������������       �                     �?4       5                 �|Y?@�IєX�?
             1@������������������������       �        	             0@������������������������       �                     �?7       f                 Ј�U@��ED���?�            0x@8       M                     @d1<+�C�?�            �v@9       @                   �)@�1iJ�?V             `@:       ;                    �?P���Q�?             4@������������������������       �                     �?<       =                     �?�}�+r��?             3@������������������������       �                     �?>       ?                    @�X�<ݺ?             2@������������������������       �                     @������������������������       �$�q-�?             *@A       H                    �?�aV����?I            @[@B       E                   �E@��|���?;             V@C       D                     �?V�a�� �?%             M@������������������������       ��+e�X�?             9@������������������������       �"pc�
�?            �@@F       G                    <@(;L]n�?             >@������������������������       ��X�<ݺ?             2@������������������������       �        	             (@I       J                    +@�ՙ/�?             5@������������������������       �                     @K       L                  xSF@�r����?
             .@������������������������       �                     @������������������������       ��<ݚ�?             "@N       [                    �?�^����?�            �m@O       T                 03�@�����H�?�            �i@P       S                 �|�=@�g�y��?'             O@Q       R                   @5@ �q�q�?             H@������������������������       �                     "@������������������������       ��7��?            �C@������������������������       �        	             ,@U       X                 0SE @P��ʹ�?]             b@V       W                 ��) @��:x���??            �X@������������������������       ����^��?>            @X@������������������������       �                      @Y       Z                    �?�nkK�?             G@������������������������       � 	��p�?             =@������������������������       �                     1@\       a                    $@д>��C�?             =@]       ^                     @����X�?             ,@������������������������       �                     @_       `                    @�C��2(�?	             &@������������������������       �                     @������������������������       �      �?              @b       c                 �|�;@��S�ۿ?
             .@������������������������       �                      @d       e                 X��A@؇���X�?             @������������������������       �      �?             @������������������������       �                     @g       n                    �?�eP*L��?             6@h       m                    �?�	j*D�?             *@i       l                    �?X�<ݚ�?             "@j       k                   �5@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     @o       p                 �̰f@�q�q�?             "@������������������������       �                     @������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKqKK�r�  hR�B        x@      k@     �L@     �c@      @     �Z@      @     �B@      @     �@@              @      @      ;@      @      &@      �?      $@       @      �?              0@      @      @       @      @       @                      @      �?      �?              �?      �?              �?     @Q@              <@      �?     �D@              >@      �?      &@              &@      �?              I@      I@      A@     �H@      :@      F@      @      >@      �?      5@      �?      "@              (@       @      "@       @      @              @      7@      ,@      1@       @      *@              @       @      @      (@      �?      "@      @      @       @      @      @      @       @              �?      @      �?      �?              @      @      �?      @                      �?      0@      �?      0@                      �?     pt@      N@     �s@      I@     �Z@      6@      3@      �?      �?              2@      �?      �?              1@      �?      @              (@      �?      V@      5@     �R@      *@      G@      (@      3@      @      ;@      @      =@      �?      1@      �?      (@              *@       @              @      *@       @      @              @       @      j@      <@      g@      7@      N@       @      G@       @      "@             �B@       @      ,@              _@      5@      T@      3@      T@      1@               @      F@       @      ;@       @      1@              8@      @      $@      @              @      $@      �?      @              @      �?      ,@      �?       @              @      �?      @      �?      @              (@      $@      "@      @      @      @      @      @      @                      @      �?              @              @      @              @      @        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hKhKhKhG        hh hNhJ[�'hG        hNhG        h8Kh9Kh:h"h#K �r�  h%�r�  Rr�  (KK�r�  hR�C              �?r�  tr�  bhFhVhAC       r�  �r�  Rr�  hZKh[h\Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hA�C       r�  tr�  bK�r�  Rr�  }r�  (hKhfK_hgh"h#K �r�  h%�r�  Rr�  (KK_�r�  hn�B�         "                    �?*;L]n�?~           ��@                            @�G��l��?h             e@                          @O@�w���?3            @T@                          �1@������?0            �R@������������������������       �                     "@                           �?:ɨ��?*            �P@       
                    �?���h%��?(            �O@       	                 ��A@Pa�	�?            �@@������������������������       �      �?             @������������������������       �                     =@                           �?d��0u��?             >@������������������������       ��t����?             1@������������������������       ��	j*D�?             *@������������������������       �                     @������������������������       �                     @       !                    @����"�?5            �U@                           �?�)��V��?2            �T@                           -@�θ�?            �C@������������������������       �                     @                        �?�-@؇���X�?            �A@                           �?     ��?             @@������������������������       �����X�?             @������������������������       �`2U0*��?             9@                        `fv2@�q�q�?             @������������������������       �                      @������������������������       �                     �?                            �?�eP*L��?             F@                        �|Y8@���Q��?             D@������������������������       �                     @                        X�I@X�<ݚ�?             B@������������������������       �և���X�?            �A@������������������������       �                     �?������������������������       �                     @������������������������       �                     @#       D                    �?l~X���?            {@$       1                 03S$@�X���?U            �`@%       *                 ��@��+7��?             7@&       )                 pff@�q�q�?             @'       (                 �|�9@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @+       0                    @�t����?
             1@,       /                 @3�@      �?	             0@-       .                 �?�@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@������������������������       �                     �?2       7                    @�G�.o�?G            @[@3       6                    �?r�q��?             @4       5                     @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @8       =                     @r�{o43�?C            �Y@9       :                     �?���Hx�?.             R@������������������������       �                     1@;       <                    �?X�;�^o�?!            �K@������������������������       ��#-���?            �A@������������������������       �z�G�z�?             4@>       A                 ���1@�g�y��?             ?@?       @                    �?@4և���?	             ,@������������������������       �ףp=
�?             $@������������������������       �                     @B       C                    �?�t����?             1@������������������������       �                      @������������������������       ��r����?             .@E       R                    �?z�G�z�?�            �r@F       O                 ��4U@g�eX�?�            �q@G       N                    �?�㙢�c�?�            @q@H       K                    �?�$Z����?�            �p@I       J                    �?,j���s�?�            �l@������������������������       � ��(��?�            @l@������������������������       �                     @L       M                     �?z�G�z�?             D@������������������������       �                     @������������������������       �r٣����?            �@@������������������������       �                     @P       Q                    �?      �?             @������������������������       �                     @������������������������       �                     �?S       ^                    @�G�z��?             4@T       Y                 pf�C@     ��?             0@U       V                    @�z�G��?             $@������������������������       �                     @W       X                 03C7@      �?             @������������������������       �                     �?������������������������       �                     @Z       [                 ��R@�q�q�?             @������������������������       �                     @\       ]                    '@�q�q�?             @������������������������       �                     �?������������������������       �      �?              @������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KK_KK�r�  hR�B�       �v@     `m@      T@      V@      :@     �K@      4@     �K@              "@      4@      G@      4@     �E@      �?      @@      �?      @              =@      3@      &@      .@       @      @      "@              @      @              K@     �@@      I@     �@@      >@      "@              @      >@      @      =@      @      @       @      8@      �?      �?       @               @      �?              4@      8@      0@      8@              @      0@      4@      .@      4@      �?              @              @             �q@     `b@     �F@     �U@      1@      @       @      @       @      �?              �?       @                      @      .@       @      .@      �?      @      �?      @                      �?      "@                      �?      <@     @T@      @      �?       @      �?              �?       @              @              7@      T@      @     @P@              1@      @      H@      @      @@      @      0@      0@      .@      �?      *@      �?      "@              @      .@       @       @              *@       @      n@      N@     �l@     �I@     �l@      H@     �k@      H@     �g@      D@     @g@      D@      @              @@       @      @              9@       @      @              �?      @              @      �?              &@      "@      @      "@      @      @              @      @      �?              �?      @              @       @      @              �?       @              �?      �?      �?      @        r�  tr�  bubhhubehhub.