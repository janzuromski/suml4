�csklearn.ensemble._forest
RandomForestClassifier
q )�q}q(X   base_estimatorqcsklearn.tree._classes
DecisionTreeClassifier
q)�q}q(X	   criterionqX   giniqX   splitterq	X   bestq
X	   max_depthqNX   min_samples_splitqKX   min_samples_leafqKX   min_weight_fraction_leafqG        X   max_featuresqNX   max_leaf_nodesqNX   random_stateqNX   min_impurity_decreaseqG        X   class_weightqNX	   ccp_alphaqG        X   _sklearn_versionqX   1.0.2qubX   n_estimatorsqKX   estimator_paramsq(hhhhhhhhhhtqX	   bootstrapq�X	   oob_scoreq�X   n_jobsqNhNX   verboseqK X
   warm_startq�hNX   max_samplesqNhhhKhKhKhG        hX   autoq hNhG        hG        X   feature_names_in_q!cnumpy.core.multiarray
_reconstruct
q"cnumpy
ndarray
q#K �q$Cbq%�q&Rq'(KK�q(cnumpy
dtype
q)X   O8q*���q+Rq,(KX   |q-NNNJ����J����K?tq.b�]q/(X   objawyq0X   wiekq1X   choroby_wspq2X   wzrostq3X   lekiq4etq5bX   n_features_in_q6KX
   n_outputs_q7KX   classes_q8h"h#K �q9h%�q:Rq;(KK�q<h)X   i8q=���q>Rq?(KX   <q@NNNJ����J����K tqAb�C               qBtqCbX
   n_classes_qDKX   base_estimator_qEhX   estimators_qF]qG(h)�qH}qI(hhh	h
hKhKhKhG        hh hNhJ�L\OhG        hNhG        h6Kh7Kh8h"h#K �qJh%�qKRqL(KK�qMh)X   f8qN���qORqP(Kh@NNNJ����J����K tqQb�C              �?qRtqSbhDcnumpy.core.multiarray
scalar
qTh?C       qU�qVRqWX   max_features_qXKX   tree_qYcsklearn.tree._tree
Tree
qZKh"h#K �q[h%�q\Rq](KK�q^h?�C       q_tq`bK�qaRqb}qc(hKX
   node_countqdK#X   nodesqeh"h#K �qfh%�qgRqh(KK#�qih)X   V56qj���qkRql(Kh-N(X
   left_childqmX   right_childqnX   featureqoX	   thresholdqpX   impurityqqX   n_node_samplesqrX   weighted_n_node_samplesqstqt}qu(hmh)X   i8qv���qwRqx(Kh@NNNJ����J����K tqybK �qzhnhxK�q{hohxK�q|hphPK�q}hqhPK �q~hrhxK(�qhshPK0�q�uK8KKtq�b�B�                            pg@z�):���?&             I@                           @���!pc�?            �@@                          �E@R���Q�?             4@                           0@���Q��?             @������������������������       �                     �?                          �?@      �?             @������������������������       �                     �?������������������������       ��q�q�?             @	       
                     @��S�ۿ?             .@������������������������       �        	             *@                           I@      �?              @������������������������       �                     �?������������������������       �                     �?                           @��
ц��?             *@                           �?�eP*L��?	             &@                          �E@և���X�?             @                          0f@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @                            @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @                          �@@@�0�!��?             1@������������������������       �                     @       "                    @���!pc�?             &@       !                    @և���X�?             @                         y�H@�q�q�?             @������������������������       �                     @                             @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @q�tq�bX   valuesq�h"h#K �q�h%�q�Rq�(KK#KK�q�hP�B0        ;@      7@      8@      "@      1@      @      @       @      �?               @       @              �?       @      �?      ,@      �?      *@              �?      �?      �?                      �?      @      @      @      @      @      @      �?      @              @      �?              @              �?      @              @      �?               @              @      ,@              @      @       @      @      @       @      @              @       @      �?       @                      �?      �?                      @q�tq�bubhhubh)�q�}q�(hhh	h
hKhKhKhG        hh hNhJ��qhG        hNhG        h6Kh7Kh8h"h#K �q�h%�q�Rq�(KK�q�hP�C              �?q�tq�bhDhTh?C       q��q�Rq�hXKhYhZKh"h#K �q�h%�q�Rq�(KK�q�h?�C       q�tq�bK�q�Rq�}q�(hKhdKheh"h#K �q�h%�q�Rq�(KK�q�hl�Bx                              �?�q�����?!             I@������������������������       �        
             *@                           6@^H���+�?            �B@                          �f@z�G�z�?             @������������������������       �                     �?������������������������       �                     @                         �%g@     ��?             @@                           @X�<ݚ�?             "@	       
                    @      �?              @������������������������       �                     @                          �K@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?                            @�㙢�c�?             7@                            @      �?	             0@                           @�8��8��?             (@������������������������       �                      @                          �g@      �?             @������������������������       �                     @������������������������       �                     �?                          0h@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @q�tq�bh�h"h#K �q�h%�q�Rq�(KKKK�q�hP�B�        :@      8@      *@              *@      8@      @      �?              �?      @              "@      7@      @      @      @      @      @              �?      @              @      �?                      �?      @      3@      @      (@      �?      &@               @      �?      @              @      �?              @      �?      @                      �?              @q�tq�bubhhubh)�q�}q�(hhh	h
hKhKhKhG        hh hNhJ��qhG        hNhG        h6Kh7Kh8h"h#K �q�h%�q�Rq�(KK�q�hP�C              �?q�tq�bhDhTh?C       q��q�Rq�hXKhYhZKh"h#K �q�h%�q�Rq�(KK�q�h?�C       q�tq�bK�q�Rq�}q�(hKhdKheh"h#K �q�h%�q�Rq�(KK�q�hl�B�                            �h@��H�}�?#             I@                          �E@���X�K�?             �F@                            @      �?             0@       	                    6@���Q��?             .@                           0@z�G�z�?             @������������������������       �                     �?                            @      �?             @������������������������       �                     �?������������������������       �                     @
                           C@z�G�z�?             $@                          �@@�q�q�?             @                          �;@z�G�z�?             @������������������������       �                     �?������������������������       �      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?                            @ܷ��?��?             =@                         y�H@�nkK�?             7@                            �?�����H�?             "@                           �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �        
             ,@                          �e@�q�q�?             @������������������������       �                     @                          �H@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @q�tq�bh�h"h#K �q�h%�q�Rq�(KKKK�q�hP�B�        @@      2@      @@      *@      @      $@      @      "@      @      �?      �?              @      �?              �?      @               @       @       @      @      �?      @              �?      �?      @      �?                      @              �?      :@      @      6@      �?       @      �?      @      �?      @                      �?      @              ,@              @       @      @              �?       @      �?                       @              @q�tq�bubhhubh)�q�}q�(hhh	h
hKhKhKhG        hh hNhJ s'8hG        hNhG        h6Kh7Kh8h"h#K �q�h%�q�Rq�(KK�q�hP�C              �?q�tq�bhDhTh?C       qӆq�Rq�hXKhYhZKh"h#K �q�h%�q�Rq�(KK�q�h?�C       q�tq�bK�q�Rq�}q�(hKhdKheh"h#K �q�h%�q�Rq�(KK�q�hl�B�                            pg@Fx$(�?             I@                            �?д>��C�?             =@������������������������       �                     &@                           @�E��ӭ�?             2@                          �e@������?
             1@                            @և���X�?             @       
                    �?�q�q�?             @       	                   �5@���Q��?             @������������������������       �                     �?������������������������       �      �?             @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@������������������������       �                     �?                          �h@�q�q�?             5@                           N@��S���?             .@                           @�q�q�?             (@                            @X�<ݚ�?             "@������������������������       �                      @                           �?����X�?             @                          �g@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @q�tq�bh�h"h#K �q�h%�q�Rq�(KKKK�q�hP�B�        ?@      3@      8@      @      &@              *@      @      *@      @      @      @       @      @       @      @      �?              �?      @              �?      �?              $@                      �?      @      ,@      @       @      @       @      @      @       @               @      @      �?      @              @      �?              �?                      @      @                      @q�tq�bubhhubh)�q�}q�(hhh	h
hKhKhKhG        hh hNhJ�� }hG        hNhG        h6Kh7Kh8h"h#K �q�h%�q�Rq�(KK�q�hP�C              �?q�tq�bhDhTh?C       q�q�Rq�hXKhYhZKh"h#K �q�h%�q�Rq�(KK�q�h?�C       q�tq�bK�q�Rq�}q�(hKhdKheh"h#K �q�h%�r   Rr  (KK�r  hl�B�                            �g@`�Q��?              I@                          �d@$G$n��?            �B@������������������������       �                     @       	                     @     ��?             @@                          �E@$�q-�?             :@                           @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     7@
                          �d@      �?             @������������������������       �                     �?                           @���Q��?             @                           @      �?             @������������������������       �                     �?                          0f@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?                           6@8�Z$���?	             *@������������������������       �                      @������������������������       �                     &@r  tr  bh�h"h#K �r  h%�r  Rr  (KKKK�r  hP�BP        A@      0@      @@      @      @              ;@      @      8@       @      �?       @               @      �?              7@              @      @              �?      @       @      @      �?      �?               @      �?       @                      �?              �?       @      &@       @                      &@r	  tr
  bubhhubh)�r  }r  (hhh	h
hKhKhKhG        hh hNhJ]o@bhG        hNhG        h6Kh7Kh8h"h#K �r  h%�r  Rr  (KK�r  hP�C              �?r  tr  bhDhTh?C       r  �r  Rr  hXKhYhZKh"h#K �r  h%�r  Rr  (KK�r  h?�C       r  tr  bK�r  Rr  }r  (hKhdKheh"h#K �r  h%�r   Rr!  (KK�r"  hl�B�                            pg@ �o_��?!             I@                            �?@4և���?             <@������������������������       �                     .@                          �;@8�Z$���?
             *@������������������������       �                     �?                          �d@�8��8��?	             (@������������������������       �                     �?������������������������       �                     &@	                           @�eP*L��?             6@
                           �?     ��?             0@                          �h@�q�q�?             @������������������������       �                      @������������������������       �                     �?                          �g@�θ�?	             *@                            @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@                          �g@r�q��?             @������������������������       �                     �?������������������������       �                     @r#  tr$  bh�h"h#K �r%  h%�r&  Rr'  (KKKK�r(  hP�BP        B@      ,@      :@       @      .@              &@       @              �?      &@      �?              �?      &@              $@      (@      @      &@       @      �?       @                      �?      @      $@      @      �?      @                      �?              "@      @      �?              �?      @        r)  tr*  bubhhubh)�r+  }r,  (hhh	h
hKhKhKhG        hh hNhJOfMhG        hNhG        h6Kh7Kh8h"h#K �r-  h%�r.  Rr/  (KK�r0  hP�C              �?r1  tr2  bhDhTh?C       r3  �r4  Rr5  hXKhYhZKh"h#K �r6  h%�r7  Rr8  (KK�r9  h?�C       r:  tr;  bK�r<  Rr=  }r>  (hKhdK#heh"h#K �r?  h%�r@  RrA  (KK#�rB  hl�B�                              �?� �	��?$             I@                           �?     ��?             0@������������������������       �                     @                           @�q�q�?             "@                           g@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @	       "                    @�ʻ����?             A@
                           �?l��[B��?             =@                           h@      �?              @                            @؇���X�?             @                           �?      �?             @                         yJ@@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?                           �?և���X�?             5@������������������������       �                     @                           �?�q�q�?             2@                            @r�q��?             (@                          `h@؇���X�?             @������������������������       ��q�q�?             @������������������������       �                     @                           N@z�G�z�?             @������������������������       �      �?              @������������������������       �                     @                         �%g@�q�q�?             @������������������������       �                     @        !                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @rC  trD  bh�h"h#K �rE  h%�rF  RrG  (KK#KK�rH  hP�B0        <@      6@      *@      @      @              @      @      �?      @      �?                      @      @              .@      3@      .@      ,@      @       @      @      �?      @      �?      �?      �?              �?      �?               @              @                      �?      "@      (@      @              @      (@       @      $@      �?      @      �?       @              @      �?      @      �?      �?              @      @       @      @              �?       @               @      �?                      @rI  trJ  bubhhubh)�rK  }rL  (hhh	h
hKhKhKhG        hh hNhJ��whG        hNhG        h6Kh7Kh8h"h#K �rM  h%�rN  RrO  (KK�rP  hP�C              �?rQ  trR  bhDhTh?C       rS  �rT  RrU  hXKhYhZKh"h#K �rV  h%�rW  RrX  (KK�rY  h?�C       rZ  tr[  bK�r\  Rr]  }r^  (hKhdKheh"h#K �r_  h%�r`  Rra  (KK�rb  hl�B�                            pg@`�Q��?"             I@                          0f@��hJ,�?             A@                            @�X�<ݺ?             2@������������������������       �        	             ,@                          �K@      �?             @������������������������       �                     �?������������������������       �                     @       	                    �?      �?
             0@������������������������       �                     @
                           @X�<ݚ�?             "@                          �H@և���X�?             @                           @      �?             @������������������������       �                     �?                          �E@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @                           �?     ��?             0@                         y�H@���Q��?             @                          �h@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @                            �?"pc�
�?	             &@������������������������       �                     �?                           @ףp=
�?             $@������������������������       �                     @                          �g@�q�q�?             @������������������������       �                      @������������������������       �                     �?rc  trd  bh�h"h#K �re  h%�rf  Rrg  (KKKK�rh  hP�B�        A@      0@      =@      @      1@      �?      ,@              @      �?              �?      @              (@      @      @              @      @      @      @      @      �?      �?               @      �?              �?       @                      @       @              @      &@      @       @      �?       @      �?                       @       @               @      "@      �?              �?      "@              @      �?       @               @      �?        ri  trj  bubhhubh)�rk  }rl  (hhh	h
hKhKhKhG        hh hNhJP�=hG        hNhG        h6Kh7Kh8h"h#K �rm  h%�rn  Rro  (KK�rp  hP�C              �?rq  trr  bhDhTh?C       rs  �rt  Rru  hXKhYhZKh"h#K �rv  h%�rw  Rrx  (KK�ry  h?�C       rz  tr{  bK�r|  Rr}  }r~  (hKhdKheh"h#K �r  h%�r�  Rr�  (KK�r�  hl�B�                              �?� �	��?             I@������������������������       �                     *@                           @�Gi����?            �B@                            @j���� �?             1@                          `d@և���X�?             @������������������������       �                      @       
                    �?z�G�z�?             @       	                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                          @K@�z�G��?             $@������������������������       �                      @                            @      �?              @������������������������       �                     @                           @      �?             @                          0f@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                          �g@      �?
             4@                          �N@r�q��?	             2@                           �?      �?             0@������������������������       �                     @                           �?ףp=
�?             $@                          �@@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKKK�r�  hP�B�        <@      6@      *@              .@      6@      $@      @      @      @       @              �?      @      �?      �?              �?      �?                      @      @      @       @              @      @      @              �?      @      �?      �?      �?                      �?               @      @      .@      @      .@      �?      .@              @      �?      "@      �?      @              @      �?                      @       @               @        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hKhKhKhG        hh hNhJ�"hG        hNhG        h6Kh7Kh8h"h#K �r�  h%�r�  Rr�  (KK�r�  hP�C              �?r�  tr�  bhDhTh?C       r�  �r�  Rr�  hXKhYhZKh"h#K �r�  h%�r�  Rr�  (KK�r�  h?�C       r�  tr�  bK�r�  Rr�  }r�  (hKhdKheh"h#K �r�  h%�r�  Rr�  (KK�r�  hl�B�                              @���H.�?"             I@                          �h@�	j*D�?            �C@                           @4�2%ޑ�?            �A@                          �E@��S�ۿ?             .@                          �B@      �?             @������������������������       �                      @������������������������       �      �?              @������������������������       �                     &@	                          �e@��Q��?             4@
                          �d@      �?             @                          �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                         y�H@      �?             0@                           6@���Q��?             $@������������������������       �                     @                          �g@�q�q�?             @������������������������       �                     @������������������������       ��q�q�?             @������������������������       �                     @������������������������       �                     @                           O@"pc�
�?             &@������������������������       �                      @                           g@�q�q�?             @������������������������       �                      @������������������������       �                     �?r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKKK�r�  hP�B�        =@      5@      ;@      (@      ;@       @      ,@      �?      @      �?       @              �?      �?      &@              *@      @      �?      @      �?      �?              �?      �?                       @      (@      @      @      @      @               @      @              @       @      �?      @                      @       @      "@               @       @      �?       @                      �?r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hKhKhKhG        hh hNhJ���7hG        hNhG        h6Kh7Kh8h"h#K �r�  h%�r�  Rr�  (KK�r�  hP�C              �?r�  tr�  bhDhTh?C       r�  �r�  Rr�  hXKhYhZKh"h#K �r�  h%�r�  Rr�  (KK�r�  h?�C       r�  tr�  bK�r�  Rr�  }r�  (hKhdKheh"h#K �r�  h%�r�  Rr�  (KK�r�  hl�B(                            �d@� �	��?             I@������������������������       �                     &@                          �h@��Zy�?            �C@                           @�'�=z��?            �@@                          �E@`�Q��?             9@                            @�q�q�?
             (@       
                    �?      �?	             $@       	                   �;@X�<ݚ�?             "@������������������������       �      �?             @������������������������       ����Q��?             @������������������������       �                     �?������������������������       �                      @                         �%g@$�q-�?
             *@������������������������       �                     @                            @؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKKK�r�  hP�B0        <@      6@      &@              1@      6@      1@      0@      1@       @      @      @      @      @      @      @      �?      @      @       @      �?                       @      (@      �?      @              @      �?      @                      �?               @              @r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hKhKhKhG        hh hNhJf��"hG        hNhG        h6Kh7Kh8h"h#K �r�  h%�r�  Rr�  (KK�r�  hP�C              �?r�  tr�  bhDhTh?C       r�  �r�  Rr�  hXKhYhZKh"h#K �r�  h%�r�  Rr�  (KK�r�  h?�C       r�  tr�  bK�r�  Rr�  }r�  (hKhdKheh"h#K �r�  h%�r�  Rr�  (KK�r�  hl�B                              �?z�):���?             I@                            @�r����?             .@                           �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     "@                          �E@���Q��?            �A@       	                   Pd@؇���X�?
             ,@������������������������       �                     �?
                            @$�q-�?	             *@                           6@ףp=
�?             $@                            @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @                          0f@և���X�?             5@������������������������       �                      @                            @�	j*D�?	             *@                          �h@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKKK�r�  hP�Bp        ;@      7@      *@       @      @       @      @                       @      "@              ,@      5@       @      (@      �?              �?      (@      �?      "@      �?      �?              �?      �?                       @              @      (@      "@       @              @      "@      @      �?      @                      �?               @r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hKhKhKhG        hh hNhJ��nqhG        hNhG        h6Kh7Kh8h"h#K �r�  h%�r�  Rr�  (KK�r�  hP�C              �?r�  tr�  bhDhTh?C       r�  �r�  Rr�  hXKhYhZKh"h#K �r�  h%�r�  Rr�  (KK�r�  h?�C       r�  tr�  bK�r�  Rr�  }r�  (hKhdKheh"h#K �r�  h%�r   Rr  (KK�r  hl�Bx                             @z�G�z�?             I@                          Ph@ȵHPS!�?             :@       
                     @HP�s��?             9@       	                    �? �q�q�?             8@                            @�����H�?             "@                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     .@������������������������       �                     �?������������������������       �                     �?                            �?�q�q�?             8@������������������������       �                     (@                          �d@�q�q�?
             (@������������������������       �                      @                            @�z�G��?             $@                          �1@      �?              @������������������������       �                     �?                           �?����X�?             @������������������������       �                     �?                          pg@�q�q�?             @������������������������       ��q�q�?             @������������������������       �                     @������������������������       �                      @r  tr  bh�h"h#K �r  h%�r  Rr  (KKKK�r  hP�B�        D@      $@      7@      @      7@       @      7@      �?       @      �?       @      �?              �?       @              @              .@                      �?              �?      1@      @      (@              @      @       @              @      @      @      @      �?               @      @              �?       @      @       @      �?              @               @r	  tr
  bubhhubh)�r  }r  (hhh	h
hKhKhKhG        hh hNhJM�%hG        hNhG        h6Kh7Kh8h"h#K �r  h%�r  Rr  (KK�r  hP�C              �?r  tr  bhDhTh?C       r  �r  Rr  hXKhYhZKh"h#K �r  h%�r  Rr  (KK�r  h?�C       r  tr  bK�r  Rr  }r  (hKhdKheh"h#K �r  h%�r   Rr!  (KK�r"  hl�B�                           �%g@Fx$(�?             I@                          �B@HP�s��?             9@                           0@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     6@                            �?`�Q��?             9@������������������������       �                     @	                           �?�GN�z�?             6@
                            @z�G�z�?             @������������������������       �                     �?������������������������       �                     @                          �g@�IєX�?
             1@������������������������       �                     *@                          `h@      �?             @������������������������       �                     �?������������������������       �                     @r#  tr$  bh�h"h#K �r%  h%�r&  Rr'  (KKKK�r(  hP�B        ?@      3@      7@       @      �?       @      �?                       @      6@               @      1@      @              @      1@      @      �?              �?      @              �?      0@              *@      �?      @      �?                      @r)  tr*  bubhhubh)�r+  }r,  (hhh	h
hKhKhKhG        hh hNhJ3�hG        hNhG        h6Kh7Kh8h"h#K �r-  h%�r.  Rr/  (KK�r0  hP�C              �?r1  tr2  bhDhTh?C       r3  �r4  Rr5  hXKhYhZKh"h#K �r6  h%�r7  Rr8  (KK�r9  h?�C       r:  tr;  bK�r<  Rr=  }r>  (hKhdKheh"h#K �r?  h%�r@  RrA  (KK�rB  hl�B                            �E@�q�����?              I@                            @���y4F�?             3@                           @������?
             1@                           0@      �?              @������������������������       �                     �?������������������������       �                     @                           �?�q�q�?             "@������������������������       �                     @	       
                   �g@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @                            @¦	^_�?             ?@                         y�H@��2(&�?             6@                          �g@���!pc�?             &@������������������������       �                      @������������������������       �                     @������������������������       �                     &@                           @�q�q�?             "@                          �P@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @rC  trD  bh�h"h#K �rE  h%�rF  RrG  (KKKK�rH  hP�Bp        :@      8@      @      .@      @      *@      �?      @      �?                      @      @      @              @      @      @              @      @                       @      6@      "@      3@      @       @      @       @                      @      &@              @      @      @      �?              �?      @                      @rI  trJ  bubhhubh)�rK  }rL  (hhh	h
hKhKhKhG        hh hNhJ	��<hG        hNhG        h6Kh7Kh8h"h#K �rM  h%�rN  RrO  (KK�rP  hP�C              �?rQ  trR  bhDhTh?C       rS  �rT  RrU  hXKhYhZKh"h#K �rV  h%�rW  RrX  (KK�rY  h?�C       rZ  tr[  bK�r\  Rr]  }r^  (hKhdKheh"h#K �r_  h%�r`  Rra  (KK�rb  hl�BX                            �E@z�):���?#             I@                           �?�LQ�1	�?             7@                          �:@�eP*L��?             &@                           0@z�G�z�?             @������������������������       �                      @                          �f@�q�q�?             @������������������������       �                     �?������������������������       �                      @	       
                    @�q�q�?             @������������������������       �      �?             @������������������������       �                      @                            @r�q��?             (@                          pg@�<ݚ�?             "@������������������������       �                     �?                           �?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @                            �?l��
I��?             ;@������������������������       �                     $@                          �h@��.k���?             1@                           @      �?
             (@������������������������       �                      @                           @      �?             @                          0f@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @rc  trd  bh�h"h#K �re  h%�rf  Rrg  (KKKK�rh  hP�B�        ;@      7@       @      .@      @      @      @      �?       @               @      �?              �?       @               @      @       @       @               @       @      $@       @      @      �?              �?      @              @      �?                      @      3@       @      $@              "@       @      "@      @       @              �?      @      �?      �?      �?                      �?               @              @ri  trj  bubhhubh)�rk  }rl  (hhh	h
hKhKhKhG        hh hNhJp۶hG        hNhG        h6Kh7Kh8h"h#K �rm  h%�rn  Rro  (KK�rp  hP�C              �?rq  trr  bhDhTh?C       rs  �rt  Rru  hXKhYhZKh"h#K �rv  h%�rw  Rrx  (KK�ry  h?�C       rz  tr{  bK�r|  Rr}  }r~  (hKhdKheh"h#K �r  h%�r�  Rr�  (KK�r�  hl�B                              �?      �?             I@������������������������       �                     0@                           @�������?             A@                          �E@�ՙ/�?             5@                          Pd@z�G�z�?
             .@������������������������       �                     �?                          �0@؇���X�?	             ,@������������������������       �                     �?	       
                  �uf@$�q-�?             *@������������������������       �                     @                         �5g@r�q��?             @������������������������       �                     �?������������������������       �                     @                           R@r�q��?             @������������������������       �                     @������������������������       �                     �?                           @$�q-�?             *@                           �?�����H�?             "@������������������������       �                      @                          0f@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKKK�r�  hP�Bp        9@      9@      0@              "@      9@       @      *@      @      (@      �?               @      (@      �?              �?      (@              @      �?      @      �?                      @      @      �?      @                      �?      �?      (@      �?       @               @      �?      @      �?                      @              @r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hKhKhKhG        hh hNhJp
�UhG        hNhG        h6Kh7Kh8h"h#K �r�  h%�r�  Rr�  (KK�r�  hP�C              �?r�  tr�  bhDhTh?C       r�  �r�  Rr�  hXKhYhZKh"h#K �r�  h%�r�  Rr�  (KK�r�  h?�C       r�  tr�  bK�r�  Rr�  }r�  (hKhdKheh"h#K �r�  h%�r�  Rr�  (KK�r�  hl�B�                             �?�-���?             I@                           @P���Q�?
             4@������������������������       �                     2@                            �?      �?              @������������������������       �                     �?������������������������       �                     �?       
                     �?���Q��?             >@       	                  y�H@؇���X�?             @������������������������       �                     �?������������������������       �                     @                           @
;&����?             7@                          �h@�q�q�?             2@                         �%g@z�G�z�?             .@������������������������       �                     @                          �g@      �?              @                           �?      �?             @������������������������       ��q�q�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKKK�r�  hP�BP       �B@      *@      3@      �?      2@              �?      �?      �?                      �?      2@      (@      @      �?              �?      @              (@      &@      (@      @      (@      @      @              @      @      �?      @      �?       @              �?      @                      @              @r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hKhKhKhG        hh hNhJc�#yhG        hNhG        h6Kh7Kh8h"h#K �r�  h%�r�  Rr�  (KK�r�  hP�C              �?r�  tr�  bhDhTh?C       r�  �r�  Rr�  hXKhYhZKh"h#K �r�  h%�r�  Rr�  (KK�r�  h?�C       r�  tr�  bK�r�  Rr�  }r�  (hKhdKheh"h#K �r�  h%�r�  Rr�  (KK�r�  hl�B�                            pg@�q�����?!             I@       	                   �E@¦	^_�?             ?@                           @�z�G��?             $@                         �uf@և���X�?             @                          Pd@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @
                            @�����?             5@������������������������       �                     ,@                           @����X�?             @                           @r�q��?             @                         �%g@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?                           @���y4F�?             3@                          @K@�8��8��?             (@                            @      �?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @                           h@և���X�?             @                         yJK@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKKK�r�  hP�B�        :@      8@      6@      "@      @      @      @      @      �?      @      �?                      @       @                      @      3@       @      ,@              @       @      @      �?      @      �?      @                      �?      �?                      �?      @      .@      �?      &@      �?      @      �?      �?      �?                      �?               @               @      @      @      �?      @              @      �?               @        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hKhKhKhG        hh hNhJ�fhG        hNhG        h6Kh7Kh8h"h#K �r�  h%�r�  Rr�  (KK�r�  hP�C              �?r�  tr�  bhDhTh?C       r�  �r�  Rr�  hXKhYhZKh"h#K �r�  h%�r�  Rr�  (KK�r�  h?�C       r�  tr�  bK�r�  Rr�  }r�  (hKhdKheh"h#K �r�  h%�r�  Rr�  (KK�r�  hl�B�                            pg@� �	��?             I@                          �@@V�a�� �?             =@                          `d@z�G�z�?             @������������������������       �                     �?������������������������       �                     @                           �?�8��8��?             8@������������������������       �                     &@       	                   �d@8�Z$���?             *@������������������������       �                     �?
                            @�8��8��?             (@������������������������       �                     "@                           O@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �?���N8�?             5@������������������������       �                     @                           @�IєX�?	             1@������������������������       �                     .@                          �@@      �?              @������������������������       �                     �?������������������������       �                     �?r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKKK�r�  hP�BP        <@      6@      7@      @      �?      @      �?                      @      6@       @      &@              &@       @              �?      &@      �?      "@               @      �?              �?       @              @      0@      @              �?      0@              .@      �?      �?              �?      �?        r�  tr�  bubhhubehhub.